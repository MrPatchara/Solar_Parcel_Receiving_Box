PK   MP�X��Gq	  kN     cirkitFile.jsonŜKo�8���Bs�V��`�Ї�i���C�Dw��Y��6��/)Kv���t32�U�R�c�X��{֖��z^mZ7���m�Ygw g�S��_��߲Y�ܬ��f��-������������j��y�v�n�+gk�]�jgsQ��K+d�+��uY�ڙ9���/)c	�VF����+W�ۺ�����R��Y�^�q��3ef��9���3G�0��5G�03N�j�$ϙ���jQ�6�k	\
ƹR��9efR�����.i�j�Fh	|���E�-�|Q�6WKˬf�6%���\���<2脝�'��03N�p6�����#M��ԧ�I���>�RW4�i֣�M���bG����<��(���[ �Dr��.�Ej�$��Dt��5���C"H�{�~�O2�f�i�'���3.#�J�_0��e+�'��Ğ���'�Vx��\:ɐ`E�����Ċ�Y�Kn	V�-_b+��э����tl%|��b�V0����Mvc��VT+7ٍ��X�i�Koz!���_�^tݜ4C�!Đ�bLC1&��i(�4c�4�i(�4c�1����C�����Q��{��rE,ЯZ�.��V���I��$VD+2��Ċ�e%�@�[��Kt�N��Ɨ��F�t+7ٍ.��Vn�]�ӭ�$Vl����^H�/��� i�4C�!Đ�bLC1&��i(�4c�1Ř�bLC1��_S�������������Y��i�v��*+W�}��ik�fw���O(u�����Ο�9�^�T�3GV�Z�2����G�Z�i���W��K �{'�6��$�P^u�`��tȤV˶~i�������r��[/MMm|�����Ew@N��h��.�'��;<7G�$?77�qt�dNl�P����b�d�.I\t��%qk�7����	E�������E_������[*?d �A�2��8�2V|����J�b	T.�
&R�Drj���T0���J"RID*�H%w$��eŦ���%tL�	%c��IL�rP���'�!�H�	:��8�f����3�2���I�d!C�� A���40h`����A���}x��e��B��g4��q�[H�>��Y��2�5t^^�ޒ�u��Kg�k8���M���>�~���U�p���9�ٿ\��@�9e���0��C|��Cb!ە��|Ѻ�^l�6�������v��7=�����+�w���޷�g�v�)3<���6]���}.������1�/l���d��;��`�KY���e�[�l�kD&�KUe�\�s���,�ɺ+���PTʞe���Vʝ���s�ݴ���\�BΔ|���\�([�W�BC�+���>t/u����A��C};@>(\i��LpSX-,�:0ui��\���r��=��ye��B��3��[SL`���H�Bd�,�����~ 
eAH�;`��4���Xxb����� ��CZ���53��\���9��D���jpG�B�Q�V]���Ձ�iw�3�R�g�0��volƍ-@Z��N
� ��`�p�G�pf�E�\#�&:�*�X�/1�K�̵B�X^VFi]ɲ�EDT�A��Ÿ^z8|��k���~$A��^��g��'����h�j�A�(9���D�S��<\X�.�-��UTu�yN�%f��I��
詁7��a#��a�ioe���#�W�k8��8��Y �p����/���{j�؁y��{�qO&�^�_�0�8����PR��a0n�q��ק��%G�DА!WaTÀ
�� �/0Dއ
Ը�g>w	��Γc�ø������#(;a�"u*`v�acX��u�� cZ;�A�g�1�z(v�j��D {�'8��/\�nvܯ'X0D���}�|
�0��8� ��%<A�@8�ܯ�g�����[9%6��u��ͳ�@4��e喾��r��)���)�����Ǜ'�||
�>Q�G:h���~{m=/���տ�����o6�˿��C���!��$���=�oQ=d���'��{߬����O�ezcn]_5w��M��)]����λ�M��ޗ�So����C��?������m���ۻ���CȜ�0A`vI����s��L��>V��'�������1A���R���Ē�~����=�:����bp��?!v��A�?�\��L��ͼH��:Q�5 �	z�k���7tT-�}%v��c1��ŎN\�R�g�i4v�~�D#.�ĵ���\����G�|�c��ߟ�e����J��_�Ky�QQXD6��tT,oq�`��:71��y,��⒏Ǧ�H��[��Pj7�����εM��n e�����տ��r���ӻ�}�>��g��sm7�qU���Vm�<���PK   W��X�Rr5�  5 /   images/01f582cd-60d2-4b90-a97d-c02e30bcefa9.png�gXSY�6@���c!��cE&�;l���ҕ�*EzO�(�t,�����
J�*5Ajh	5��Cq�yH��~|��o�./=g��ֺ�{����g�_����)�	����9}Bc��`�>q������ ��f��W]`0�S�o���a�=�3'�/yƎ�pe�00ٿ�ڴ��E�=��͏;����1SV6�[��`���9��w~�K�*�%�6׈�Ǚ#Q#�˿�Mi~?���u�Y}��!�+�~"|P���%�1[�ߊ{��}�z�|�/�?�X�~W�@z�3f����jC�?m����q�9���?h�lĻ�;x{/��YBS�"f�uF����C�<���p_�y'7|ÝWj��x���3M��#t�R��s����W&�j�0�pKb`��/{\y�T������;�g^u/��*Z�~��n��M��JH �h{�;*"�t9d
9\�fMϚ�ċ��#��.�]'o�&&E�F���MܓꝨ������8�➣�ϟ��X�g>�1��W"b�������9��p��ut"���xx�+w���ȳ��!S�|��r,�����ʫ��Fp&���B���R���!F�$�}��K���!��N�����ӷ�U�$^f*�=;�	��n�X�w��r�ܟ�@ԅ�kW��O�ީA9���D'ԋ/����W�}�H]���ǉ�3�P"n���t��j8��ܕ�l���eȔ�ћ����=��L�6b�E�h%9���Þ��3w{������1�I-�v��,?�+&Fp�g��؊z
?|��AT���{v���!�*%����زkAf��ΛsK�f��*���-��O=�BRO���'�^�Iy�y��_�1K�/�6����`nkk��1�	���Έ�8��8		��U$�1�hk��v6�M���9׆�<TI�歈4���ѹnNZRQQ�v��V�k}�T�ӥ����،����y��+��:B�JO4�4d
]\PX~m��v���ޗ�W<2w��@ʯ��E�3tJ]b��3 <BnDv�L���QVA�*?��mV��oߜ�ܤ��7iL֗��bV�������O>�A� ����ۋg�����C(�����[�I-���
�a��=[��������=FVfO������l�R�e�F����2�^l|��W��\ �N��KOx+��M|�������C�Z��n�G�������-9�C`>�:ឰ[��q�a #;�233���C�s+��0���?��M�^�VV�ec�>��
)��sޥBR��.���8�Ԥ;�����魶y�9hu����<���=)�r}�ֆL��J���M�ܹ���3�����|)����3!�1�Qi&3#cpk���C�,B��`��!Khǫ�W��\�|�}=D'D���~�i���R2�H�r��"�Qc��D ��W)Y��O	�8O��$�8Drqq:C`P>싄T��c� �H���C���J�֬��zhxh�9����Ǥ��J�$Y���t��"|�]}���A����XoI�� QG*m�^'f�;�e��/V��2��у���
^(+I�|ǿ[*�\�	�)�<l"�����x%�*���,���Xߊ^�(����}�L�'o"�M�n��[1!U�����n��*>�eQ�U�o�-C�e�K�t5:Ӵ�3R��n-�.,�+�{X�ݐ����Xh��!i��-mH�G�9�q{#���s�K_���G �+��oQR� y�P<Y�4<<��<d�2��N�ݩ1rS$�wcfg]'<J�޽��q���鷅�s���(AQ���ǰ���q�X��/�ÇoR���UmV�zh�2L�6�iF
�`[��}�f�}"�d	�@w#������}w��&s�u��?E�]�����!�Jg#XU����48�Ю��o]��~m�"C�8���o�>����f��M+�#>~~�����J��n�j6H���#�hP��F����[��|<Mo~ u��;1�Z�����r�㵮�H�C��Q�J�zb�O��4\qr
b̥6���@����[�?�U���ë���[���i��S�����C�D�W�I-��]*�ADS��q-����ܛ���ɱ�3�4
�P�F@y�o��f��i���q��*�痨i���ϟ?�	���rV{�6��b�/�A�\��&����
6�J�[�)�<tOH���t_�n���t!Js��H��;AiD�*ixk�C6!y��ґ��j;�H�A���C�i�WIt�B���h;�+�W�#�#��<�;U%�^پ}�p�������KM���������l�M�gS���/���@jR��뮃tE���rvl9��Ձ�;w�<2���J�Z������} �I8�}���a���Jp�Uapz�y�S
�YgK���]Y;�I���U!�~� $��b�������$~u"��L�(�QM���@*^ �@%�|���VO�E�{q�K�&q�peUU�.1+�eH��ׯ�S[^�A����4a0��Ѷ�3Isss��I�����n�U��L��dû�O�K`
0�[~��Ͻ������Z\����3�J�C��ի߄cy^�a���5hp�v/$�һ���o1����3>~S̽4Kv�kHK��<����u�*��K{A��#U�,q�A��F�p_��/_�<b��)��yqG���l*7��!S9�|�3��M�Syyy��١�6y�Z�l�aY-p�9��(�c�Pu/P���a����o���:>�Y)5��+�����Ӭwi����{Q��7'v��:+
�`��e��I����h;���q���bR���ה8��h�8��Zx�2#;�@{VR�|L�TJ���ϰ��;�`����/�,(ƓwNӅe���.�������zw'��F�@�]����&�п�E��K��bYk�m�=o$~�v����Z���|	̙_4(l��]P�gzf(�5O��]sp�<A��_+޿`y��mb[�Ļ@�H������1?�Y��xC�T�8I�{����j���V|jii��"p�Am-����`�73�e�M�5Gr�k��)װC�(q�AZ(���IF��X?�����ڦ���ߛ�znF��|�T�jm)/݅(��oPRk�ǹR�)��-�.�m.�N[��0
����3�}�3��SS�S���sR������������Ġ��x...�q|暰|�m���b��� i�@�ZE�$��T\�}m&�յ~`�/��؎��[K��HB�����6I)O����[a� �fW�9X֥��?�K-�0��(voKB�C�fa�R�¢"�Q����X4-��/�AFs&d������Oi,N�����q0vA�[S�A7@��������p����T�Յ�'>��<�%����	�5G����@�^��簠�Ck��R�ხ{qϩ/�&��ri��A��A����o��Z��A�����e���t��U�Ty7}]"�d���%E�S$�%�� ��ڦ2{ %pC��y��d�ɓt��x�q .��L0�sw���>�I��ܥ!��2���s_�{����Z���!y
��c��d��v�TO!�(#�?~���q�ѭI�[�6�L�ي��x�[�2���fп�)�y��(|*ۼohx8�A�{k��B�H�3 ���ݢ��^>mJ-���n*�O�����!	u �&�8�ꪑQ�nkF3�Oy��bV��|���w)��]!$^W��_�ے�x�Sm�����ʈw:h[�q��-�d���4�c�ǌ+��XI>v6 s�>	��S�!��,?��B��'� 'ȴ�@W�3����?¨W�"ˎ-a3�6^��i/��+M��O ߟ�,��^��A`�&@{�d���]/��*$�����z$D<*y��Y�]ւӭH(qy#�)8'M�`&s�,��s8����ȐY�?텽�cz�@�T�'�PO?�N���da肝��Ŵ����SS]t�L���,�_u�ЏԳ����e������rM��f�!"����L�~dd�{��ٱ�լ�N- �gK�Ր�$v?|���ݔߤJmVUn�9���T�j٘	�7�n���c��~�[x=�����P���0{�g\�niS{$<�e��|Vv0~L�����Q���]^ᯥ��:�Ra�T��5��2x�"n���9�LU�cuʦ�eQR��(��?�J]ȗ8B��Q��]mZe�nVQ�F��ֺNj7�c�!��,$�4��H��ߕ�0òw�2{&�)	Ԏ�`��T�J7D��������A���(���G��HH��f�ڙ�/*DxvԘ� 7G���B`�w�^ñ#��ުQ�QȞ1S�=Ȇ��.������t�t����|���)��2��݈� ��8�8oEi!ߞ�q~c��g����:�EJl�}���~I
w{���٬����F5�E�T���ʐ:8dԬW*�c�j���j{�3��'��M�j`�cY!e`��|��L����y��ל���Z��U���VnOCc�:��p~����4hֳV�@��{��Mf��& :��h�Ε��B║a������O#x<��O�w���TZ�������p(yf�l�P�X϶��`���A�3U�I ��:NX;���W�k���f�̓��Ntip��(�/��<���S-(�
��>`�N����R\xo��US�T_���d����FPd<�-��zA������e�Dv�O�N>�/���iS����O?�aV[
�Oŗ��DY��Y�_6�1���O�<�E��ւ��ؠ2�[���4ogI�ߖW3Q4U�O�;�-�����b�t��Hp��r��Q3RQ�3
�]9虙�%Z��*p��3�B��S�
��@����!aaR�q�0K�&_��f�׳}��|!V�K��M���1�K��!�HR�VL�f��̯�(&�ίS�eJG����JFNJ�R'=x\U��M<n$�9��ms��N��N<ם��S$�Rh-aI��xb[���:�+�� �za�����ê��*���i�ղ�x-f��w��t��MX�$�`�L�Թ*?�(wJ�,R���s;$�e�qr������
Y�^�s��Y����G�=�]"���2e�]�j��������z��.��@��p�l&��SC����q�
M���V�g��I��� �^�E��jF����#[aV�*Z^�l��8��v&}�I��	�� Z&p�f��L�\��̖��7m�h^O5Ͱ�Ɨ���M�Sq�G���Ŭ� y:4�ߘ���En7�������FIkf�l�<������\�;�Bv]��[������G7|^���J`g�.	K�ӟD��8q�x���T�-��w+:��-+K̊��D �J�J�|��0�@ufP�,�?ڈO(\�,��Zȧ�c�gT��ʖ��^��[w�a�K�{dvB��u��E�Y�O�X��\Di�:�n:w�ɗ��ʞ���֖����O��H�/���
�|y�b?��J�hp��Hh�@?����,��>ګJrQ5�7;H�w����9.'S��hs��1g�"T(�q/�Ka#�e�I�֬@��@� �ݫ���n2ȇ&A%��v��]��f~�i-ٞ?�d����x˱)����G�����D�9T�i2U��l��9�Ւ��^ \3m�4�'�7=�2��\�R^���6Z�,o�*9P���1���Hq���y�^�d3_D�'Ee�kQ��㚜�.���:��v��8�M����Vh�B��R�M)���;�U�W���u�9���]�l�=g�IɎXD/�Ӽ[Xi�"�DX����5G�\�!s��K��:@�$�fޢ�Σv`��y�!rӋl�{c��o�t�c2+1m[ޑ 'I�U-�k��6���wM����iR1�гFUI�MXC��5P��N3Q �}>/U���X4K��K��	�h��&�� ��v뢀ڲ��@�]�Y8��0)��-f�Z�V�����E#i��&g�{_�]Y��Rq�z�{l"����!�d����ʈ�~c	�i���oIO��`e�Yy2�ɪ�n7n����̳_�
?O�T��5(7��?�2��X��E�ٌ�a��]���93� oS��(���ń!)�̞��u���Cm���%V
:v���&=��%7����'y `f�1�z[j��e�}FscЛ��M}�����V\��Դ������d���˚&%f�ӑ���a䲎H��b��w.�̯�F�$�q�$�yϔuQ��b(4��C��dU"��
�b��R�����sr�q��V��7��?W'���s�ϟ�'Q��Bc�bckU��fkkCV��u��wx��XA`:���Q5����gEbM)?�"�&]¼��]]��PVmE_��i&Eh�n�"a[V���'%�/zU	yD���I�CIn�\YG����Ls	�49{Gc{h�E��2��(��n����x�����!�5���.��s{/��n���p"cϪ��͐~����C��
B���<?��~�kW�x���ny=\+�r�(zxM}s�CP:�ϛ�������KK��2��b!�O9ҏ�p-�AξQ͹��|t���j�<�tF�q ?�.q����a-�sJT������kB�͟g�}��K��A��[�3���J�
H5,����M�=J��4�$N\��L����rT�w������zj��2�)�r�/u���eg7�u�1��ng��\7�`U	'|+%[#�
aD�]W�,#���K C�;09�~k^�����>Lc��H�n���ޙj�������Q��1�EV��7	y�Hl��x�W�i$�}x��՚�$����TeÊ/��M�!K�n�:ơ���"�
���Jm��#�1�~�p�@�b��cR�X�X8��._ҡ|։Y&�% ��|k������lǄ{��};Zm���疨��YV���x%`ɘ�f��BI˞r�,��/Jξ̤TӆX���e��q"T���B��u���[��o���D���Es���~V��k�ۦ@��>���Di�����	G��bl\���j�J�[픙�
�04�I�k���~��hX���x�|�i�ϒ�V	U��Ɂ`B0Y��X���Q��h���	%3��5�w�>57E9����j��B��S�cs��0T\t�P����˪|{=D�3�LҖ��c�0vZ{�߽!>i�8QLX��s�S[0�VH�����z���?knn�E��ץ�9�;��$�o�c�I����9�5��G��xצ3yx�z��������#y�Ǿ�y�n����kQr0+\������,���=�@9�z����_��r�l�6W��2?�ӻ0	W��ߪ�3}�***��y�w`|x���Ws�������hj�æo���\�:�����A!�SLm��;,BcmF�.]��!�/p>�dԚ?�#M��S��'�T���a��(O�g%{�'�S����U^���q蹅P9TsS53����ؒ���=b+�0�n�#T�$�*U�Q����Ȯv�n��ǜ)��Kh��r���P�����ٷ,��U�4n0Q,�	"=�_����&�������Z�U�a�3���-��_�og���3! �ǻQ���x���*w�?m+��=��v��҄�R�_d���Z'�2��q��T��m0ٝ�OJ�|���\�퓇"�4!�V@�-~���8ʅ*K��v�m�:�fl�7����6�PZ��|:2
G�I�.��Jrݚ�#Z�#��H��a������i�q�N-��z��e�$X�)�r_K�W�@�"�dz੎�����?�O�>W%�n��+�WL��=��q����%���Zʻ�BY��M?��ϙ�ϯ�O��m���t`J���p4��a�*�7ә�#�ݞ�<��1>�F�ULY�<�(+�� W.G��4��񚩓i�����=L�Z��287E'�Fhow/M�صkׇ=>`z4H�
A�/k�����X��i��#��b&#�,�Ͼ��-S�������~V���}6P�U�4(�w�ﺥz��֐sZs��֗��]!�%� �rrru��+P��	To[A�����\Z=�[A�D	�b�uW���(�6�O��md֋x����lմ��a�g�� $dp!r`wS$_����P*ݔ=.��?���y�w��w=�8��O
�ɩf�w�9����|��#Z#�Iw�k����m���J�I�-D�>(9M����Ip�S^��T�irz<�A�g�� <���_eJ�ٿi+�B`2��?��{����EgQR�l(�?��I_{�#VI�Xu4?P�奙	U��,���
��x,�d�<b���K�ӡ��D���1��;|ϻ�E�|����J������N��>smF�=-P�iKjvl�ó�>���G��4�q�̏S������ts2j��{Ks��N߉μ���~��
ٚ0�7"���+��o~�΋����^^���:��=��p��pyQ����^�ޢ��,�e��0Gi�]���N��� �_��M��&LG�D�;�4�`^�P�Y������h�[8���$��tx�2���YB���ԍ��f��U��<`�xt1��$ߣ?<i?�)�Xtn.~�7^c*�;N�Ñ)��Ս#�@P5~�6�X~���h�h�3b[��i����!RH�ZPB�{����lu��T�l�^C���R��9��+s��o��hYA�`�`��
:��}5��5G���C^7��J~�ی�(�ݞ^�>Ѕ%Ш���\q_/���`
9�. ��&�Wρr+Lq��o�މCS�Ķo��j�x��*#���a˥_�M��¤���/�fef!=�C��/sI��s�G{���s�s��{#���[a]?J�.��$l�a=�o��_����afg;����P>�4�1��g�Q	�]�ʳ�����F�{�8��`gg��Oȉ�,\0���Rv���wg����K�j�!D����-α��2Q��vg'!�������g�|�Iw�]w�[����7�|v��>c���\�f������h��Oފ�Ut���gNK[%(?y}ՙ�(�9aWCs�>h4-[J{�Sm�U�}N��f\{����p����	���a��L@h��j�uT��-'�W��,�y$��*���_��.S���x�lykq���d�b�X�4�V�?�'DF���|xA���c���H{�� �:�kb�"���{�[y^��;	��zXݬ�h_H�f����?�(�+vظ?��ך���Dn|��m���b��JRrE����4���S�������A�|�Ҭ��#2����T������*+�E۫f&^��
B�XVr�m\�L�*ѿ ay6%���K�bUg{�Vqn�^��QVfT�Zs&��9z�[gU�����é��c���S�J����
jw�uJ=�-Sfjt�}��~"�M�w�0�S�r��X�r�t���U����\5]�aJ��){TY��oN�n".`�+4p7e]��!$�����0���3��$���}bm��EϪtU`vF�.Wn���9ӎV��`�;{�﯅�?P��
��^]��4x��T#�>�L�U�c]��o�w&	�G*z�A�I�B�����bWt�XO8��9�,?��*WMU�Ȓ��'߾F�z�{U�N�����A����s��۸ڹW�Y@��jy��*m���d��������YXC�d�v�Bs�r7B���:b@���}��I"��?-���Mޟz��,���ݱc[q!��󷽃��A��&K�:~�^y��0��zT��cx�&�<a�i%�+qc�.�m�-e��|<	b֕�@yDAg�
X�_~OqM��p�t�N��c?���_�����!�eW����̯_�[���lpX��n��Y� +�z7E؝U�*�V�ʷk�Lh�7��:�E�&���"x+�&b��T%U�Rbx-��Br�?�p_���K��,$�|@���1�0F�=�Χlا�y�/��Q�g��5���d*�~���O�J:�ޥ�ث��S���ga���4�#���� �J�]�*	�����gj�1e~�;���e�����P-�������NE���ϟ�"8q�Z���
q��##���F�C�y��T�8��"D���Kw�����ذ��b{��O۷9|[8s,u�[۔	�P�Vib����Z;�;?um;��B!A���=#Y�*7�0c�E�2���{��d&�&գ����Y٭l��F�<C4Ԃ�!�gt9�׻|@���K�{�|�>nZ���FZ�ު�<��M����S������HN|���S:ZZ�����J��D�m�������X��%��Zh�(-��[� �$�,L��q��a�Eno�'M�A����r%�/_�Pa�����X��,���14�z�L��_	3�
GBc�9�}�2���S���؉y䠗��/0P'��YS�y�@�΋��W�����b��qc0�*>
R�3n��S�W���%?�{�o��	�p`��|dlaa��V�Ԭ�)E��t��_]��P(-hڊr��S��7.��i^�*9�:%�2��N�"nmSn�58躻����ܺ����.&�-�Țz@�e�^Nl�=vâuv6ׄ�S���	����n�;��ϲ��I�����3����O,~�r�"�#�ڮ��N`��}�I����8�*<u�L���U7�S^�j-���9a�2�A�����si�Ж�T%�jֵW��
��������֛lWf��9�T#����%�$���za��)֊OG�\�h끌n�>�r4M���W�׻5�c�l��u[���w>�}-����=(GX¤O�������W��ڜ������<�S��ڌ|���Z�����#�B#o�e������v�k��7S��|]XȂ�%�,R2H��r�@��^[���l�� T�����n���b��U�y�7����O�q�
�׷�+q��aD�w��^��C�w-�	��9�X��§4�����s6L�&v����[Aj�u0�w�eV	��ʆ�.��X0d8/FV��,�<��L��E�.w}�ڜ,f�k�!fM1�_�܃�2��Ҋ�fQ��t�5��d�ن�s2��.T�5M
4�m� �6�RP��Ջ{��llR����ŗ>n��� ��;���f���-�1��K������|�y1�(�����z�31�S���1b}��|�@�����V`���ֺ��`�KG�o�@(�X�F�I�U�Y�)F��F<��`BX�j.Xq��>�B��f��=�<��Ԋ�_@����i�L�uK��6���p�]ߝs��՛��7�x��i�!'�RjJx��%����Zg�2&��.g������VffZ���}lBB��_oaw�4�^xg�Tb��Eh�I���E�Ů&���cZ���C�i��\��+R��+��p�����h�����i�}�J�Z��C~a�D�����R�N��A�����Χ4�=,,,:������]^���1e����D�v�ι����=�α���%�����`;�=��V��5C�V�m�oo�Wi��ko�f%CW� `�P�B�r(���I�o�a�ݿ>g�"0|�s��d��Fd[W���V.m/�]�wh4Rt��R�����A��ެ�r��l�߯�U3-a	�'�B����RSS���������}��uQ�^���cc&���ס�4 .�.Y֝w�����(X�!���L�5�����Ֆنd��w]
 ��?��f���,t���R ��}=/+�Ɖ3#��I	����k/����q�Y���Vݜ�5��X�D�RN��|g����|�_�'k���1K�F0�zi)���i�ӻ����J��xv�eO��M���[ <�S���!�M�ϸ�f��)�M�����=+oy�}�$���9#���γ,^�]ap3�1�ݔQ&�t�q�_>�: 6%L%f��<#�c U���\��`#��CkA�lV�x̲8��%7������"�/��mϦ%�հ������}�.���\� 0d3����'?tp�%P�hk�=��7[K�S���,��O�R��RpO�
����� ��˥�|~9X���;;��$�����R9H���z�{@;B�\����<���P�up�O� _�,��v�Sܻ�&��5��LL�fH�n�� \#�)���y#��n�@���gIY�z1��|I_���ye�h�}(ZǾ�w����y˯#D��H#E�A�&�%z�k��''�l�2歐2�	��&���-8ǒ�Jg��Kc�~a�c5
�o1k�7���!����%��?js�*�n�����I/[āMD#��۷?]y��~Lk�D��q7Z�R��$q�׷Ma�@pM@��U�����!���xJ�~���,��;j���:�����PM��MS8k� ����ۅV��Y��x8qm��E*FN� �(d� p�h��vG4�P���J��S�Rq���yUx���UV��Y0�r�`�~�5>h�\L� �~��� �1��5H�A���h��J�P[��\����L�B��3�+4ӱg�o�+���d\hKt`I���~q�z�u55�e��-��8�J �����:V"���?ȍA&��2�v��i/6��Mh�E�pU ��_9��do�i�Un<�n��	��؈� n��*����V�L<�B�G���NǗ�=��[��v��Պ�!;���p�:�Pٟ�P(x�l��K�7<�����i�
0���:�֞�}�{���h�7G_�l�Hg��?�dE��Ç��6o;��qs�k%�Uj��Jom}~�-�]ɱ��69%ki���º��Ɵ�.z1�(�_Uç���>�F�Z�W�#��T�G�UXqa�Ǩ�����͠�r=�8FxT"YZZ
�n������?&������Y=�A��	9��던��:�ʬ��/ �:�q߰�5;ui��g���5w�����&��UI���w|�"�n�&u?|��,���)++KV��5��v��g�{+�(��a��[�M��r����I�_���CP����M��|��"�3UC!�$v�^i�5��7.v�(�SI�c<�����$���rb�A��w7Re5`hi�`|1��O��V^�pl\��Õs)�n@R���:��<��B�QD�̪K�?mt�G�k�oq���65��C�vJ6p���+�x :;8+[mr��C�3P$<B�_	��r�MD�Jha39a/C �[�b���
敞�$�*@�v�nn��bC�}�������s����8�Ř���<Z��q�R�]݃�� E��脘A��d1æ�G������8�W�U9В��vv(���Q�@RI/d�w����>m���Mp�$��֦0�_e�1�Yx�jk)=r�ު���[�J#�Bk��ur?�Ņ�Y=IT�'�`C7�s�]||U���[u�hk�T��ֆ�g�c"���Zn"���[�0`j�/2Z+_��uE8�fx�&+@H��d'��u��M�y�����8#�z�N��SM���'�L��E���0_ ��Q�3I;���Ҟ]�ګ���,���U�χ�T�V��ŋ9V7�s�W-4���w>��	���L�Nq���-�1*�k��614x�B@*z�hY�`;�j �砉�4� �Y4��U"����NtHKéu�o��i"�?v0RCr1��)q�{�ެѱ�b��.���2%U�3�0�#��f����5M.���S� �v�}�.Ũ_��_�E���B���� �W�h,͛U#;t�xW�> '���nD���V.���jj���_�EQJ>|���ʜ�
(��|\v��2H�'�2�PV�0&�f`KO3��s�K綗����A^����_CϦ�N>�Ry��>-[m��nݚ2��Qz�	��/��E|",��:T�	���}(�|q�$}��f��U����aЁ�<��	��gϞ�F���1��,d{� P�ak����B�`/�8�"��o��������:V�� h�d<Њ~���8�zl�"�ZLh0�e�Mo����{ȈW EDGE-����������>}�F��J��E0[�ѐ��w�tGH���)[K�i=��p;
J�~6���#A<Zɱ!��~��6��Br�fC����G��<Zꘓ��@�?�͐)#F�7g����S�r��� Lʒ2�r2P�	I8n�����N5�E�O�%
���D(�=#sm��%h��O���ww>!�9�Jg�h<�9�YU��Q����-����m�>pW���,M�bt2)�����T�AVV$��I"���H��y�� �����~'�NWd~\B-����A
c�.p��onbԤJ`˯�6��ʮT��`�ʊ����nm�׽ks;r�Uc�wQȝ��eQ�R�^� �a��@mZ�Ǐ22 ���f�4%�����9���s.Dg,�IjW=�498B��|gy��/gv����}�%$iuׄĻw�@Ƽc���O��#�v�*¹w|�)���O8�|�2**���^���� ��9L2	����s�'ԗb�[������L ��t���m�Ɋ[�;~S��E�h���!�}�����JY�Pk�z�/����Y[D)g8��t�0jJ���a���B�<��#9�]�~�2���q��G��U�gQN��~���I
P����V�s��=�h�b`��Z-�*��'�)�0p暫��;1��P���gc&w�����k�������p��Y9<�g��ۆ�i$ZOo%�� ٩:))	�a��(���;�Èn6~��C_m����Nw��Y��8�����!�&��]�G$$d��F>�cM�pd{��^F�W����5�zԞ�cd�>̞Ԁ�y1�e���P���Ǐ�N�ǭ՜@�3@�R(���|5r�W\96�����>��;g@�����b���z��.Z�����!�J#hR���^:1i��ō����kA$g׫H��YD6�
��p�D��=*�ZD^��N'�0�ݲ[�`�_�Ɂ����6o%wtt@ (j{�����KX�{ 1�f�V&_�hG���ȩ�m�]�~�c�0[�Mr���������Z��r��i���_��vHLc���/|!z�1��+�1!R�S�1�M�
x�`q��<�������h���j��l���uQ@+:�ʛf|Ĺs�V��������[��ϝ@U��:�YP�M�m�������P�pR	����C��*�%?�m���AKG��0N|-�;8wlHj�[8q�mm2��� 	JII�mLUKL�l�al�>6"(ʹ��M���\�`h�Q���-��C@+1̀����.f���)KM���:P;0�e � *}I2����9`��n����xP��Y�\��:r�c���	���.��<9��M�
���0��얕��cW���՝s gmሥ���6���-���� 1���V"�/�mY���_�Í@�&�w<U��ܳ�/���b�3c{"a�7n$��Crઐ����tƞ��'+��1������O�lW�v���q�P54G�CƁz�B�>��1����a�o"�m��,��
�BJ�N�Z��JS���|�T<Dֆ�:�'$<�μ�{7tl�wz\Mۅ�Nw������5cD�J�Jb�62� `�f�ՠ���J�*�2��R��m�f��Ӷ:)�2.��s�	�D�=� �OA�?PO�6ܰE�I	�O�t�f���w<F����e�e=J{�`	��2�geiY=7�V��{��V����SV��y�ӌY�_�|95���5�4���{3��x�N�6���!�#5j{@%ܭ�³!)����5u^��wE�~�+_��������C�9��9}��J�(�z�S�����q���*�j�W���\�#X�;��˿�l}w?4�}� A�nSt>5">{#Ѻz+y,�xr�����,ݏQR�KHDf�C~������n������n�-y���F�&�����ˮ%�����daR��ųsO@�	���\���_�8_4A��0L����!ن����E�����? e�=�{b#�=X������P!���ǰ��,��I�ٿ]��XT�fgg?�T�<��a�ʠ� �.}Y�r�6��R[������CI �z�^=/=�������h��$���߭첲x?�#�ːWz�lT�,���y^v��(���\���SyI��9�ak�-�4W5���G,d@����Es��'�y�ůQ��ړ��@��p�N�&w�~.-�=a��.ʊ�&`&.u�쇈f�+���(�?~��U�Y�t�@;IF�����UǾ�e��I8�L�Hܦӈ����n.55�p���oXƀZ����2�:��܌
p�=W��o���I����𫃱܁	3sm��X���IVsgY��cS�R72g���j0� �O�p�]��ҫ�]XRR�g�iQT0Fc�����Hmmm�3dee�v���+`ԓ���쾬���|O`�"�"��^ۼ�/����LJ�v1o\�����������ԕ�'|� Uo3]�¯�@��ެY�.+˥�E �lލ}w���	�[��}�&��+����/�ۀ������I�=s��K��%f���<op˵k}$��>2��+C��v�c����i�BKY��R����>��	�9����8N�F5��8�?Ź�(6Ѭ�$x ���˱�
�>�XˣtJ?|��7�����J�^)Ֆ �ĉ���G�1������CI54��	q�������������B���o%�8�,T
:�S^@�t|f���8��w(V��Q��D\my �9�R��ح������k�OX����hK5���Β?1j�l�j]&��Kr�0�����v���ZĊQ���'4��8��=t�����2�L�ؼ�ƂN�tڤ5ϫ��o�{,f}�~�LW�Z˩G�:Tol�q�w*��+��tm�ݓ�Qۛ�������Sǜ�n;������|�ϯ�"�|������5) �gP�|�C�F�ǳ�V��Ro	�pDso�L���ZaR��!�ύ��P�/�_0�=�-�'�MY{z�|h�7�
��J[v;o�b=z�n��|`僉I�^�-������$�Z��A+�g��12t:G&�ƿx�@!϶U�v23�:�e��-Ӆn�'�l�l����jR/k�� �G�Yv�uX�w��<L��[�+�j�vT;��Pw׫܀%�Lv�B %X����ɏ6�	�`۱��r�����㡉����Wr�o@NV��~޲��|9��|I�u��Kw��rͅk!؁y�@�;�D�9qO��x�]_О���ej�>��^�f��Ce�Y��uZ�Y�N�z�~ {�1��D�!�m��OT�:�0�-�O}�:��`�*+�](���
�ﾔU{�a|�t���:�w����)g�oD������U(Z�5Q�����Ui��)?��G��k�~� !`;Q���F�K��d&�YAb�Ԗ��ă8Q���_�MD�2�X�}�՗�4`6{�ܤ�{x�A� �x�fkи��K_�fW5��'�_tI�y��i?�p�J�?ҁ=wJܺi�7ϳ�[sz2P,�U	`*a�@���	�8�<�pb�e颃������+�/�й���ZS�G�^�z�vb^�t�_��`߼���eq�ѳ+�/ج6��,�@����p����}���"a>�I5/�X��W���M�;�}��Y�1I���1�Ţ�vp>�7O<�Ϧ��1�ژi0��z���?��G���������c�l�/��G�����S��vڟ�⎯����Q��������9d���D^;�J�������|������<�o�kZ&�������_�/��K7�6B)�A[�/h讠����@�P���}��g�J- �^�B�6~͜�P�X�`9C�i���q3p��'þ�	e&�xb��2�߱37�p�Qt����كI�Џh�?e�j���Mm���ل���I_<�`�3saoV�h�e{�ɼ��]-O-W�����հ�0	ߝeb���vU	_>�]�2��8YL��:Z�G�gD�w'�� �c�o<�G�`a�u�xV���n�cYhe��s��r�:ߕ�|t3�וo:���U�wa���d~o�-���.ly���gWT��z.ݷ���6%��Lɇ|o��°)*3���Gc�iP9װ��#S	�2���V&QJ���Ut��kv`�[�����2ye����
�>q�>frYn3a�7���ٵgΖ$�sjM�)��2�u�늹����bK���yE�Y�-M*��^�*-�����k�/w����G���?_\�j��W�9�+#�k^s�:��K�Ŏ������#�]o��wP�e�����x����H��H�
]��u�k�|���#(�2N3 ��0�������Ҡ�����L��{�x���oܒ�rJ%���J5e��TR)�b�(��3�E%�i�u*E*[�)�mB�uƖ���e�>�g�,Α~�����������i�������z_�}���G���)��d���$10h���|�мM��v��9A!��Q�i���(V�7�^��ϣvYN�<��mڸ	!��s��4�.�	E�\<�dA��^H8�o�%�$P;۾Џ�OP��2L_�Oh.L���DJ{��c-���m)�+��f�)l���\�/k=��&P�P�W_aV��F~��K_�N(��´P�˸7�A����&)Y����6 �(��ͫ ��H�}��
ӹm2,�Y��9��H�}M`E ?TeZ(b��h������J�s)H�������p�b��X:p1�b�S˯\8��w��"	`�&ȸ2�q˧�o��P���Q�7�!�
�jQ�B����J?��B�N���ݤ�ϖ&�����X��/D[��y����:��ꍖ� �,�҇);%��%8`�;�����g�>}I�`�'9����N�ǀT���C�|�%��i2��@2m��3�ˎ S�f���&��G�B�	]I���k���mOd���S��3>�~��b�5���oTo�^8%S-����Ya�ԫ����D(2�~�
`������7���@I�G�Y�6}��`%��V*Ӟ�h>�(�=��P�N1�	_�A�ΐ����g�,L��]`��S��s|򣊸yH�eqA ���S;��~!�a�����29��0k�Zim�Ef���S�4 ��%����%~ZP$�b��T`��~5VZ�o�O|Ԏ��*0hC   ��ڝS̾�`q��hq�{K;���~�wp~�wp�o�'i�_�|�w����������������������������������������������������{��m
���s%�k�~Y���5�?���HCW!E���p�Q^4B6��������uGV~�@Q[<kUf�4G�3��s��6��iD�O~}�B���C�VJ7�H�bx��+P6�Sc#��C9�ъ(̋�Lg�t�h��FЇײ��^�����J�ݏa��\�Ջ�I$K�������TJg8��� ��=]9rY��^��x�@��N6���2Dxh����t�bΡ��v��xy�I�"Ngxe3��z�57�ч���>V��q���_?�41.����M��o�_���DD]V�tȶ���m$R_#c��¿l}bA �Y:���,�k��5���7��S��mo��(���5J��Y�U9�yb�*JR2�͜�,�p�~����س�dϽ�L�`��;HV�)L���SD=L�)u�\z���Ǯ�La_�H��%�ӑ�TZ��|)UPĥ�6w	��wiQ2.w���f|��X���$;��^��p�z�h'�?Xjϴ���D|�	�j�~~m��pL�a>���jė>�{��d��]3� ��|�6ᐇUX�2�9������-ԑD�S.��&c�B�43��GOM��̡w9�y��.P�p_�2)v�~��rťe���1�h����S��_<�߸�B�	��zǇ�rG�́�m�Xť��TN�E��q��D�$��R;��<2������	y���]7���K+m��# ~�5Ц�����%��>��[f�[w]W��~6k�s�O��n:S0_=�����N�2;'�˲�\���a�5��Hx|6��3��;+OmN�B�s yu>X�.1'j�]^|�ΰޯ,��8�����4�<�s�c�nw��(�ۺ�t� ���H���>-�4�L�sZ�I^������m�u�v��y�4���үc��^��x�na7g�sr8��T�w���������#5U:#vS�q�v��fAL���J�	� ���#6HN���m��ə�ϫNڕ�6��<}�mO;�_�����"���W���ե��h�p��٬�i�N0K��Oy�U(^
ao��h���k�|���T��ې-Kt���r����u���M��iYa���Æ�v�����X�Y����jrS�W��7̦��<

_���_�s��D�Y͆w ͜Μ���K�&S�!��۸L�{�i�����L�a��]���;V���	sl�=��4�u�9��Qng��2�����6�X�ι6�~
9Z?��j�ŚAt*�����6"���J��0XQ�c��'����������"���c�]gƻHb��ױo5O���o�5h�I�OIh�0*�����ϡ-<�~��	��2�o7t�$�nz��P�����EȊ��Lu����S#=�a{�j����L.1x%�J�����cǸ�z�j��>���1n���>p�&�UGU�~)�s���ʄ�u�Hq��M�@8����w��7uk1Z[ʵ��818 FY彌2��s�������j.�"u[[ͦA�%.�+�G@�;�+^���)������"O��рI��3\x=,��~5u��t�*DW�ϑ�=/��t�(�]����E׳��CJ�'�׃�c}L��ȿ"��3��ׇ����<�ZVH�ͪv_HvjŎ�*����I��Tck�}�� R��H��"7�qe`��x��S-�?�$:�a�Y������橫_�X�1ӶZ�g�OA�� ���9=�b}�Ž����ӿ��8~3`L�>�[A�0��e,���렞n���4�|C`��7.c�����4gNU.����b�V@5���%��?8�!S��$�@�D����~�Z��������^[P�$���Ϗ�o�w�G�ȫ�7�\~lԥ����/3�"|E�(�����K��@=� �׆�u�����=3�3'(��BE��)�d�m�S 6$�Ћ�M)# ����v�G�	_���:3��<_	q1k�_��8��P���#���S0���z��:J�j#�P�f�]$��r�ـ���ˡܠRfTZ'�_Dz�'v_��?�+���o�o̎��9�<*�˰/�B�uʸ���t:�H�V�i�FZR~p.hi��k�d�9�[����e�EA�ňA�p*\s���ݰ5�|�V5�J��K�|�8����"��#��B�Ǜ���a�4BsGoP�����"��_J�vm�@���N^-ř������<<T��}|�*˂^�@�9���vA>��ee�r�ELtF�fN|���Q& ��:��,�ǿ�DA~S ���Q�+��iw�ŉ���9�s}Į9%	s��]<l���� �B�E��/��$��*�q�-�9��a�� �ĥ��?T�@Wd&�����-�z!����X�chҙڄz�E�5@Ĥ�}p��ȋR����@
w�b�`웒�j�e�17�S��4��p��wegHF-f����*�@��o 5��@���`�*�o˻~x�n��5d�]�/d�.���i�X��ߣ���"
���jIWM;��K�O\ ���k*�T�K�sj:�p�,�%1v0R!�\�h��c�%��!�-�(mW�o��?A_SHṞ]���)�٥�/:>G�RP����rۆ6��=:|���x�U뵽h�jʫ��d��R4��ޗ�r��w�d4����Rr�;�zqQ�h���ה���T���Y5V��g&�=���qB�)��)|�i�j��8�Z�У���I�j �G�k/��v��ig6H��`�"3J��<��s�z݂��K���Ik�Z�I-=��,����]�!�����íq���`Y��F��Y�z}�ǽ���m�8O�gX�y�k���wf٠�=�II�,?�3
X\��˹�����H��$;tȰR^�vט�7!bbF�m=����囲�x@=o�	b#f�s�/+/ۖ����YC���E�w@�-"�*D��IǍ�і�>����6���qc7���Y���}�	�m��9���)���(D�5T��ܿ��6(�sT.�yB���ΩjY��~���#ƙ��Wp_5Yb��O��x�bL�������m�v7y)�; -�E���t��=��bEE{hi�
�]hDl�c%@��
D��1p��>����;cđ�M}��H}��'OL��~���AtGp���. ��w��{�\���)��(�b�����X���t<�������4��uF���%{�M�4�4}���>�M�:I +my��L�w_]g���f(,���ݏ�KNNb4�B��zg�a	���[�KS�/�)�
,����h��o�S�����������:w�Z�Y�ET3�n�YKl@!ˇ9��/)Z�gݺ9��\���E[�����:���"B81��AS�H�CN�vD��V��gsKqN�Rȋýge�:2��N�_����9�H�*4����Zc��$���$�69[�^h��÷a(�>�dN����O�!��"�g�a�+n�,Zn$�e_Vۦ^�v�A'�o��i��_�[z]�Tq�|�O����.U�~��z���e"��-w�}E�q*�'�J�_��2Rl�ðq�B��GU�sΒ|�$���
�a�(���iU����e���A�,�L��/<��c��ayJ"��J��/3Н�i�3T��]��8ǘ1LF��]�w��3'�H����PA�@"�ɬ���51�'֥TX:v%Kq=��ڵ-�B���$;l��&U1&�2�qx�������M���"=.���p*.]�	�bw
�$�jċڧ���<%7UqtB�;��»�@�R�츽-;KQ5T�hw1��VIy�8�-�c(F��_��2H:�Ŧ¸��dp�l�$�7"�I�W���/�d�-���^wc	(���ަ�1�n-A�^���A���o��f��!9omKC0�ӆ/�a���.F3UC���\�U���i�)ͧf�U�\�iZ����I�g�p�]��Lݼ;.����ʣ�T1�������	����4�� ��!���z�9�%�5��0/$�R*Y#-�e�����F4�BP}s��~�?5jԾ��5Y�U��M�LuOdl�&�a�*��x��O���T�:m[��j�~�J�e(=K��g�i�\P���h��z��g�d&�s�&U��hH޽E���?yaQ��P���[q�-��� (ǜ�?�������n��XzME�{u�J�ؠI9��1	�����D��>���Ɏ��NB�N-�0c��x���ƒc6�*���| ���j� w������n-P6�G���
ɣ�O��8�ml�a@i��Q����ī���^B/�)�9YG[Ǹ�;Y2��m^�ɦ�'Ҫ݃�N@ �TV�l'�'"2C��uM�Y :�m�<����3���sQӂ�r�C�<�q1�`o���0l�5��{�k�VFJ��b(�5�����[�yy��< \)�v/��'�pLǆkiDnҙ���ܳ��(j� U�ޒݓ��&��jS�q�T0�<&��nq{��΋�Ĕ��W�B���e�L/F}���,	2�Xk��v���������L�9Uw"��Δ��n�J���.g��b}�|H@X�B�Nُ&����(�u���-���;�hB��iZ�9������⥖l�/`�GU������v�����e!s��*��H�H��/Fsr����T'EF0 �*�j�;���Q^qO��ф
��ײ�"6���{�K�§���������WxA�"je ,O��Ս8q����|N3�I|1�s��l�o�2�|���v����;Ыb+];�n���;��®�;�
tl���9����{u�j{s��\�397�004�p���:#r-+6{/�ŌL]V��!�^_��Q��m~���:\�2jpR�{��Qo��L[�i; ���u�@�0�g��=�.hF�?ba����P��CuQ�.J�������g�%H�yM�@��:ř��o�/!md�p8)Q�������*3�/%��yۤh!�s�y%�/���y;sNB�㬉�<`�W���-%����� �y��F�+���z�G����@�Yo"i	�.�����
Ԕ��S$�<����/";.�rކo���ګ�{j�X�Y�1)�J���g���(��+�洭�u�'b�:L#��X������Q|��h)ë�9��Ԫ��2/,K�;Կ-H��/���%px�J����w�5��:K��'W��&��X���N��g�	������N�����):)�褫d�F ��<ɸ���`�AKE&��:ܗNNm	o��}����������.���k���r�W�R��������p�A����$�p�.��\f�Z�r��|D�w�(��'����4Ru.#5�;ʤ�Y�O�|Ǌ�:n��z+��ͅ��#��]�;G�]���Q<�qɺ3㷘��a�쥕�=łt�2����?�mݝ�	y�QZ�oa�7��7!=SB�{Y�6�]��1�N��h��ӂ���dj�s�2�,F|f��ݐq��:.�~/��z�����VP�ʹ�:#�M�_�Iu�D3�4�����3�(��:D�n��f�n��)f��!��e
�����Qǯ�-���`���8jf�50����d��t�I8�b����(����ʥ9�P�)mݮ���o9��:25�P��xT����Lk�7�nÕ��`P����'�.MOs�
y���0���P���R_H1�HD������w��^�Bby�=C�����"偒���"Zշ-�����Hsu��I�@I�/$~�PV��sؠ��m ;�B�~N�W�s/^�I�����c܊���ͥT�%E�{�ݓ�	K������.m$����+�D�%ԝ�7p�(�����e*TAG�%T�B�,Q��K��ė*��>��R=��Mä�z��p}�Uw���pk��6oi!o6���t0*|�0����72�v˻P�豑��qd
)���:w�A6�Ie8
�	��d��W�?j�&DC��=���S�D	��(6��X�����̱D�,t^IM�@�&�sq�4m]vn�$q���3��>-����%��0ﺕ(<94X
Cqؚ�*^[4�1B��?_���(�,���{��Hɮ!�`�)N [�}:�o9(�~�丨�f���j���;l\sN��Ŝ�'wʍd]�utRG��W�@e�&jw��� �o�Ȓ�p�\E(��C$���X0�%���k�.(\-�°#�d�Z��W�D��L%���|p�rH�V�׺@z�9��IC=��q��R�9ւ'�w�gC� ˢ��kϱ#4��Ӏw���R	9 ���AsK��8��~��p"��^�r~��&�G�����J*�y����c�biِ�.��6.zՀl�9���L}S��zGvG��f���㨨Y=���)�=8P;Tҳi��������f��Hk�R�#<��.��8�~;+�ь{�XdC��E�bV�I��2���=���^~�E��[`�q�.�G{��Nr�>Ms7a�6�Y�=���4Ur�f�Qn<�h>��`�!������!#�92��VI�>��u�*'�_/D��m�����A`�f
����5a���힡4cƫ�0e��;-�y��{?�B�8�҉���x2��.@�\{�������~�g������>w���\�k�9\F~�E'B�:6����T�_&d*�sZ�p�t��C
����M��!?))�;���}M��	���/�Mw����ٗwiѼ��[�1Ka�6�C����{7��ן�ߧ����>ZIH[jp|�x����p�E����ҳ,�C0wh���'�c{>}Ȼ���������m����"�sE��&��R�q@�8� �gԖ]b��+����U�x�mu��K[G	0���1�A
G��"�dA)>м^��&��Rb��(�ҭ�#l�Ad8qe�j���c����='�%�h>
�y�J�5��@�f#��̡��/m��WΏ5��ug�.�o�UC��Bԉp������Yz�Y��c�/JU�����r�u�Z�����>���x7���X��ŏ��qW��P��3��E#�4���0^g8Ҏ��Ҽct��Ls�E�)�h,��j���ewe�'>�=���?���w%�*�C�'�x%ځ{�ۛ�b̧?�b��X�DV(,����<S��zW�i�46�0�M\��o��D�>�e��33�����o�y��e2�f�W�����R���q�鐎!���M�^e:wWV,�l}{�w&������գc�{�aJ�{���VH� �)0�繯�`O��_4zNZI�?N'иi ��� Z�����!>�ɰ���:L�M������ûs�x���2�����<�1��"?�C_+�"�2\���Ow�-ǹ�0��̡���0E�V[@��ǘ��ߓ5�)�|!��У���&YT�@�X�%�-��-��d/o�*lx϶p@k�l*�e��/o �Xo���B|0w&>X�Ğ��y�b�0�#	X�����v���G�NM k�i@Й�QI֘�X�O����
��4�Qݍ�\����S�x%~"2 �C��U/�<b�Rǥ-�/�7����_%{ջjX~��3'މ��*>���/���%��mg���k'|3�k��d��(qs�H��T��縨d�e��&���T S*�����6E����j�/�� ]���������?��N-���Ŏ����-&n@�U.)4ShI�w���Q�D�+O@��
���6lQk�;y?�r�QCn�ܾ�*�����ȶE*��=�߹d�t�m������$�Ћ�G��+��x��(M��8���]�Ǯ�)E����Q�Gح��#@��_2����yY�}�RL�7x��,��q��I�yH^_z�iA�eJ�e��L���D�������>��oK^�X�Y�"\x�I�5�glEwe�ͅ��)B�]U3g�%�B:s#���|���e %,����vձ�p;�0 �T�y��@EU?������3)v��V��4�C�V�@�L�	��7�I~����奬އV��ND���fe�$
��Id��M6��[v{�2]�eH=����e�L�:a"�e��qQ)p�7
卫�>����/1��1V�Ά�Z���)�ÿ?N���k�ȶ�.$S���+�i�=|�rʜ�N��ܑ�X���f��%�O�'�y���D��e�
�c�2A�E�Ih���Rs��lM�"�����RsE�!*`Lվُ"+�����c"���aA2��==�q/����U��2n�\�{U��9?�q;�����V��������ʊ���9w�_v������ʒ�~
���{�oi�?�F�z88�E҆�	� ��q�4n�36�q�h�`�10�.?��L+����~/7M����@DD��A�����Cs�KY/����2u��@��V��'����8��J����l��"=��h,��JG��#�hȂ��/�ؖAM4�a�#�#��j�(��D9RM ��1I��$�.���1�Q?M؟^$�����o"#p~���p����u��!i$K�X�O!�RX*�=�'.�)�R��#��;84�L��`�۷x��^XaSH�Ta���DT7٭Ӧ� ItD[�~�fagط�����K+5P�e��R�-�=a<���Q�D�$��	��
kl��v?y�����y�SZ�ea�;���-�ha�v��.�x����G�#�-�4�`��y��J�n0�o�H�Ⱥ+jD���[��5��(����cc�A={A���:���HKD<N8�IͿ�,�c
�L��|!;9�����C2_i3k׵u�L�B�ք�NIe]۝�2�KYk�K!�+���7��^߆b'Y����tCfdA�!9����� C��=�	i����joGp{n���<�#��솣(Z��w�a|:`���k�~�5���%���j�Q�hn�b�mD���d����DF�f�bD���>�>����`��6�2�>��!) �Aݏ�����~J�zV37>0�4�DnyOV��<�6q0��观^l=�3��v�Md�����(�f��D��<^��pi9��Lj�w�	O_��?�}��y-�^%p�ڋT���H�G�������}�q��a7���`�NH���_��
f M��Հ&|����b�p����+}6���]Z�m�,3t�{���9��&�0��ɂ1��D.� �H���`<'�N������U�Xd����s~Ặ�2�C�� egJ/),EI��.�l.4���"9��FH	����Q�=�<�
qY��H�ߩ��<���[ۭ�kW�R�o�I�r���E�������F��k���=�q���t���0��	��7��#�#�f��x`���_
��([M��ss 0�=3����q/�;;Z��~.�� XU�|Ax�?]�G�塹��f�w2�0��ć ���A�(�&h�9�H>�x�>m�JMT1���޸vM�gH�`�J����?���BY<K�ё���ĴIÜ�m��;z���泏}L\��SI�]�Ď��FD�����o?���Ə!H^i��'�^#��=�\�����V���t��V��t���*ZH���*����*e7���e0���˴�r�?z�]��!��D��Mz��V�*��<N�^�4�9Tƥ�O.aR
��*�A�hI� �=,
#� �r������m�h�n����6Hi�����w�7��|��Ț�oonn�<�E�������z�^x��-Ýek{3��޽령Rn)K��(C�Z3��N}�u���q���_ļ���2˅�L*���b�x?�̬��#�1x�z
ű�F���b��g^}ɈZ���Q�{1��Q�ⳮ�9����N؊����Q�	GG������#���%ƿ��~���[��$��p����
�09��l���A�1m�y�o@�Y��������"����;_�-e�KL���1>��ړ� `���Z�v';F������7�����kV�A��9��PdR���`�Am��ɲNN6�Nn�����Ci�L�k�a�=t�Ui����w��=�����T�֖�-lQ %���L���A��|��Kq%r	�g�sr�NB>����K�I�DSɠ'A2��/l�w���v�6�8}�y�Fy4//O�Vw}pp��Gy�k��i	EWG�����`�F۟c_�`V�54p���`8�����8����J�'V	�E�������{��@��`䜩>�=��>�Op�\WEY��qሻ�cV�z��a��~Ŭ�2��"~[p����J]�"����x�dZ�<~��Q�o!��#��f/�,�R�҉DU�,�9*)+k�s��l�p8�>���p<�������:�杔ɗB�L%���/���!-�x-����R	."9��}}?w�NK�Q.\�����䇬���j���\�����
|�E�F����脪f��2�/��W�X����5��.=_F���c� i�=���64��٩/0ht�1�������8Y�w�ߧ����
7��z��}[F�z:�C�Ο9Ӌ\"�]~��-n��,q��fgeg���<��ݚ�X��ny��gч��蟞�=qB/vGttt�c?��0�A8q�SN^�W�}��+�KVVV~o����g��}|����zj09�Y͈L ��T��<)n���׼�u��C�>��yk������uf�`j i|a��tt?��`煍����+++�h D
_���s���G�LM�������*'2MQ�����Q���&D�=��J�9���'�Ffgee�w�V�9X���>��h����4m("藰+J^�|G�L�e�P�'�_����eP�[�U5ǚh�O���W�ÿ�,����u䘋�t���&k�ȃ�� ʖ��j��/~a8~�/V�����?HJ����M3:�|�� �����lL�Dΐ��s�?i����B�����_�ߢR�`a��2�A�v¤�b�U��V]��zig�qI�n��u]
GU���s��j�ɑ���8e��3m��u��*`�Ƕ*}f�ۛ���ɕn:d�|����9��Cr���1Z�ϟ�9��9�&d��2��7W�k�����Nt@�*��Q"���p``�/t����RcS��&��C��`�B2�d����G/.my^P�����`©����쯥�p�Z�
�R�=&zIkruPgO��֦c��H�B�����d��lȉZ+����П5�	E��rY �>��/w&B��
��� Ͻ��a1�l��S�r����	��g��W=KK^�t�DC'�����/_�{�^�Vk�J9��zȌ[�⒙P�D���v��W���x�Ģv2�k����R��;�!% �nX�Ӥ�/��_�τM��M~���mt�T]<^swy$���p�e���>�2h�.�?��j�����._:���L���^��
��bu�;lY~�������*lpM�>����\���+SI.��72{&���r��4U��+l���>�M!��.���w~m�VU�H���HHpb�e�?3�溇�,n<H�Z�����L$+��q��_����Ҳ ^a}o���H}�.�+E�_C�oY
�B���P�BavC��Wk���s���UNٯ��I����_`(�h�i z������7&:��V`w@���do�H�����慨¯�3�x�#�J�v-\��4�M��oi�Ǯ0������t�[ղ����Ė9�*Şw�{%����u����gWݩ{����Y�|BR�b����"�._I������gϞ�6\UVV�績�����[�B���������`a�Zn~�Ⱥ�a1Jf?VՍ$�]�� ����nXM��tｻ�>}b���7�H�0�k��H7i[�� o��7�2�OJ�-M���O"��o6�JO�l���S��B��TH:>KM�e��z˰�"��'0+��g�u�㷡P1`��m����k�[���B|Ѕ4��O�n�"��j� � v�����.@��7e⽓�Zi� �J���jwru΀��=���aȍ?I�\kn^�g�X���g�ee�K�w�hW=Jg菒B�Q��ل����M̉��&��{�_�����{_�*�:��TU�G��:}�g�I�n;�ߴ?W@����n�YC
&~z�a�^��:g�#�[r�/@���q^{k?E�͊�M��|��n'��^�%rU^]ũ(��t���`w�z�����n>�O�5(��@�����5�:��w�#�"5��C����L��la���-j�&3�[ FA��X+U�)�s=�*6��`�%8И��U����7�J�VΨ�}K�L��;��4s`S��@�T��y���j�@κ���yU��8qv��
�S,`��+�)�J���>�t�k�+�9����v!��SRRR���x�ۧm�s��g��6r�k���h�`��[[[S�q���N���S������}O�Be#HZ1ۜ����@ྡྷ��e{;���C��1���/�����G~��|�?�\�����8�c�̳� ���747;�S(Y$8W}\�1򐼱M���Tf�MM�н���?#3�y�4-��ׯ__P��*��s������r(���������@�Bc䪩�*����� o���9��@���5b��.��1I�Z1-Wr��'��-��Ϡ������s���QC�*�Y��UG�&�a�	N����N�y��U�Ï�{��Y<ӒY�?xz��7��S����p�Tt�����@:�k�`7+Jn`�J�a�W7W�c=�U9iͣ9́Y������{�p�C>�7���`�B!����6���X��̮��!�_���I��1���������8�8;k`���a ����m���Z*�GG��b[[�m��������|��w��SO���� �9"�FLG����s*�o�����k���GH�S�sw�x<���&3:��SY��zj���@
R�b��4ȧ�-�[��bT�Y	*����o1t���@X���=UH~�k5G��^��m��� �Z��s��\s��"q�Q
/��݁����;M��bʁ$��;�KG��|����&l)��啕������;��w���c4��nQ�r=�� �a�w����TǴ��A�"fe-��Ao�������oA���<��T|j^��W����D�x�7)��i�Z�2�>i�%?㪾�~���bm2�H'-w���V�(_wj�9���]�ozNk�~���u'\6�-1p)>�K�`b-P�j�P6$=F�=�V�/��}��ԞZ���ϟ�h�S|�~��3�:�����rR�6
8��;rqs�����{gX���G9* hm�����v��BP@Ab���ޱ���f���L!�tf�	��s#�P�x^]4�n�����+gd��g�Z_��v�K�Ә@�k�;��C�ڣ�㴳�3��tO%r6�P���xk���qq"|�1N��|����/���Z)��+ŕ_�Q�Im3bK���\Yed��L6�y�!������|�7�\)�(����nG�L�}XS!�EDFTX��R����)v;gd�_�<�������nzv6e�,�@r{d>�譓g�^] �l��(.��SI`j�����e���4���7>�8O�x�?[W��g�猩�.�h�dw���O9�ŋ�<�ܡu����x^oՌ�^��[,�e�����0#�:)imu�Hў��tB�����8�Wq�JN=:%���x��K3&��r5�6�N�R��:�s�Sp���Q��L\΅����5������wl���w3rG��6(c��W�Ő��Ҡ��*�f��6w��u�b�٠KQs�:t��.m�&�Z.+N���t"�n7��ߏ=���e���L���?���1?KI�~��O /T(���qž���ԻSR��-��7����u�=>��ΈP��G�ֹ ��L����M��S�Ug������G�&�s�,��p�x��^k�@ħe3��9�yy�#��T�4�R@Eg ݞ�ǳ��P���.��i	���$��$dFH~����s�Ң�������O����ƾ��:��0����,ZY�N��ܝ�f�p,v��]Z_�rT���
�~���?̤��F~�٣�H �����2g��bc������5���c�E�g#fL�3��6���PE->�r� �*0��3b��]����J.�����-���<-9��C�ogtg�C!1����+uoQ[̐&#�f·�B�0��j��� %�6��PǈcJS�t�ڇ.��g���U�Ote�/_0[L�YY���ba���λ����U^�_�Z=�w�!P�vB��GϨ�N�=�� h�k����퇀���,$��ܤ$p ������9b�5��k��i�a�ȑ��ܝg<!�;W�X�\P�࠸����K:a�`j���Dd�B�d�G�w@�ƶ	݈��f�����3���Q���Կ�˽��6:��V��@P�O��O�&%<��g��?{�����'�o͍�+u��}���S6e��
����n>EN]&���QŠL�9�I�YaU��75Ey��ϗ�����{�7��2��㓔��%���O��$���Г��	k&f�ӵ���Q��H��;u0�*/[���Zx�5"�J�G�\
��;lr��@����8u R�TR؀Ϛa ���Ѭl#��Ġ+�A�����8�8���1]:�CRb'^;%�$�W=?��mPJ!9MM;\\R"�m��x�tS�Ё���=��;���{Bq���M��!%�1*�n%b끹zyL�k�kr2�?"�����.��d�U���$��`�q��I�+a�w���.{Ѱc~�M���b�?5̧#Q��̾G�oke�C-:�X� 2Uo <�$��$z\�C�����D9C�J���X�AR92{�R����ѡ�9"�7	�H�'�8���T���I,�r�������:w�"���L/��q��s~�� �sv���D//���Ass����5g��JY�AZ���QU�/.yo�Z�w���&o}�.H��W�	��(�`��:j�84��
zh�������~�v���ڒk�kd¸!!R�n�|�����HVeb��6����᤯41���9Z�n��hzbj����ֵ��=�B��˓P�E�~wK2Hv�;K�2�Ν;����Y�L�*hp̺6�!�3��?����w6X	I:::�[.�R�rJ����[U�`�F(G�l�P)��p�v�zn��	�z0d�g[V���>hf���چ�;`����D�}����|�,���?L��y ���	�=� w���P#O��yQl!��Ri4���f3�n0���7�RZ����x׭j�$FVǖ�"���Ƹ.�%L�>@�_j���L�m���޸���<���_�b<�����m�������~�CW���o�o̴�x/ڒ8t�ژ��y�ڿ�YRR��^)���t�͑B2��z~S$d�ſ�IheL<��͗N��;G[|6��Y�8`~�E)Dxccc��`�����W� �aP����<u][s��%7 ��IW�k��t�� ʷˣ+mX�@)�X2����}�G
tX�����B�(@R,!N��7��9
�Sx),��
��
�����G���p\�re�-����ij )���^�w���3%$���� �{m��~∣��_e��Z�ּ��t����_�#u+(3Oz�6���r��M@RC�t��}�3 �k׀��}�o�)%�`7�{�f2�@B|Lb�N����+���d@L��u�J Z�����H8ܭ�}L@}��`y{��]ףj�u�Ha��w�����B�	�j���ڵ�Z�;�c��٦`��O���R.Z��D�E&ޖ�6�:�%��͜��1�_6)�n[�7�A��Q����t���I�.���?�}c�.����%'�^�-U`L�.���2\ ���um�m�][��j���|I<���)����У��v�u�F>�W�){A�{�X	 M���f4	bȹ�����v�'>���؍�� >k6�w>d�H5ǚ���z`̪�LR�[�uSyyy{�x>t6� ��4��tE����[u��х�,uEbm���D���а���.�I�y��iruz\*t���[gee]3<�����fg�X�����Ii�ZqS�P���O<���A䵁]F���lN���dm�V��1�����AT(� �W?���=V�̗���Lr���Y��&�3���~߫�R���]�֐'�i�f_. �L��9�1%k�����WE�)���umdWN|�!wz�C�B<F�f�4��y�ھ�~S�l9L2�J�&���Wa�RT�X+�Q2p�T��q�o<@;f�X��+�cR�C��C��" [ؗ�VF�@�)���.�h��$I�r0�*Ր�#ץ��m�I����]?�#]F���:e�2�>�G�,a������w*.�,�lVY?�yXl��I��A�r���*7��L�%����<�*JJ��:*-�2�5&��jdzU���jO����33����gö�$[i\@@DԪ�����a�zVo2�~C$P'yxhBڥ�|�e�$���g��K�z�g�xi���_ _�3�T����rg�jE�WPaT�N��%$%!G���O���J��贿�"�wK��nH$,j�W4-i�Xʋao7tS�ww����O��_n�\�~��R�=�������[~e:�Z� 
�	u�����?L<f��V�I� ��y�V�ؐl�ȥ�:r�z�J]Ʋ�?�V|h#.X�L�����*cf�@Ĝ5���z@@`��������$a�=�K��O����^d]еY%�,�!Ց��`��?�-���k�cÞ]�H�p��4Q�MM�6W����a5=Ыe���ސl&�lhmݔ��w�%[�p��u�)Ӣ��2V�H�c&�v����u��06p�����um���!���@�&�|�y�bZ���x����s�+�җ��
זoh�{��f����^�аu�n݃@�\p�/��%n�>z4}�n~h[��Ͼ�j��a'[���\�%75�Ng��юYO$�`ۏ�	��$��2�)�F� �����\Ⱥ6o���l�����Z���*Q�zSӪfn^> gt�j��5mh+�t�e��hր�rؗTu!ҳ�VX�ݺ����H�v_�C<(d����-I�z������Pb1�i�wD�w���k{���)
�HLJ�oooO�ص('p�����5������݇$CK�v���܀�`$���SO���zx�f�i��\G��Kg��*�e2���4_]�B�ބ��V �߉�xJr�Xj���1G¡��� �_ޟ6k-e�iw�?0A�1������V�<� X�27�.��,��5���^��i��{�R
�-ҳ�]��}�H\	�E���!�g$�����;R���)��E_�迄5��oJc�ϖ� gJjA6T4e�����wU��n�Og��ʾ��8
H.�k�%�Tx���������{i�_}\[PSG.8�ibe"1�2�f�L%��A����`)H��%T1H�S�1�!� �(�$r��J����#��B`����n��I���y�Ӟ������'��u/X�k�jbgQHA�/{�;�����?k��·kt��GQte��b�o�j��u���m���h��p�J�.ݰF7�n�=�+Dt-,z�����Գ�Q��ϋ��<B�M�'��0��t�9Y�[�' �F���r�ɿ=��V�����~¥B�r��"u��6����%�p���x�4[�0Mۄ����F�7����B�_��G�dx!���īZG&l�A>(�5�DB��� 0t?�\�ݬ�e�_c�' "�� ��f�B�;]L���ڜ!gr���9�]{j�R_8qHHHD&L�!��FV0lf��G��ܸ+P�)E������nvE/�w�v�f+?Y�9�Qs�$O�|8�i�Qx�m,�U�����ϗ%�;�������@����N'�Sͪ��&㈮z��7�	�?�S/��1��_L�4�|�L�:%���'�ʇ�m����������$�l�\��D���.)|Mܠ��C���َw �{�y���h@��'�ۯ,KV�W�ZW�������xR��~�1���� ��2`Z%@�kX��Sخ	�V�P	���:�޾�}w��9�ьA���Bp��	Ϧ ���Qg	�KsZ��T�\�V$�-����nQ�~,&wF�rJӻ�p�䋐ƐK��Xn�k>=k���7�UGWvT��{�3��BT�*'��}�؅�Sw�߽$>_�o7����������8b%ؽ��>�][]�z���2� Tu(
\ݖb�tZ�ݾx}Y���x�T��K��V'Gmu�@ݥ�{�Auʹ�_�<�3�9�!��p�a�t�V�)v~��W�������[u�C���[�T���j���!��NA��կ�>�w��Ĳe2{���Fظ���c���PP�����k�+�܃m����C_�7�a��v�Zss�;U[��N��S�)����`���HR#0S��;Qv��U��of��C�f�jS��q[o�3W�Z�O�A{��y0lPA�q���j�����9��ּ����Tl�`�GMx3)�"�	�L���DՆ�3�7��^�n	<�CUF��Ff����G��-�w�`A�Y� ���*�D�y6d�N?й6O�T�g���\�o?�QbS����.V@����Z�o>�����<z�ǣ��fs�Q�e��lAϗyr�F"-p�qUTA�T�;z6��!+��^E�٥"�U�x�	mIq� i��Is����.~��Ħ��`)��u���'d�d�H�|�git�Fbh���"��t�?���b`�	�A!��5�~Ĩx��|���f�L�Υ@%���P�aq�D�0�=eB���2���8������QSc����d��b'W=d�Z��x"#�y5���PK   8��X�bZ�b �f /   images/32499b6f-cadd-4b9b-b4f1-e31be966db26.png��T[]�.�P܊C��/�]Z�h����8���+�.��)P�).-A�	�����s����ތ��+s�9ך�w�|TQz��I�	  p�d�� �'   ��q�k�������� ����Lz�K  Y�k�j)�4�س�AL��<��b�Ʀ�� sKk��.����{EvEG)s+kY/g�w^J�^��f4b� a�G��� {;A��|<�3�����V�F�� -E���$���j����{<����`q�sr��y��<�����<<�?h�9�Y�I�����3+WWGA0��ݝ͝��l	� �s�99Y)X]<\�=X\^�� m�b�l��jq �976�������]���?l\��O�;�0vs�������C���l�/�f�`s;s{sW�GZ�h� �+����?_�7��(*�Ϻ���C��*����vQ�t4���@ܜM�e><����tGA)gscW��:b��R*uq�q��[;�A�]���s�ǗͣոY�9X9��9���\�������Tbfm���G��)����H}������Hlf*hq�7~\�����9������6
JA� Ώ��p���������������������� ;�	�+��?+/;�1��� �)�'������S�?��;���r����ch��?��p��$k��h,���;s��Y����Ʀ�[���_V2���������|w+s�����A��pu7v6��|\��ѝ��ʃ�s��u���%f�=&���MA�'�$1s���������� HƲr������5�G��T��vd����)�����wo���"@xh/S�_�_>{v��<<%q���E�FM�	�K�����=NTH���^�w]*^�����ݩh�/��e�(�2�/f��&���5�5�nǒՉ��b��u���h������̠ ��6��'.���$�@����;^𿌴���E>�����8�᳛�6l�L1�N���|�FG΢��gk�"���M��k�Nm�P����HY�7T8��&������A�����7W��jH�������]|�8%��6��Pj���m����n��^x��Z]{]t��;���;N߁�zm,0P��7
������+�0��21j>*h����=()>~YY��8�Ι@x��2����y	�ҧ�I^����xԖ�NRѠ��L-_M�a�%WF�-��~��_3o��h�w��(b�ʩjh��n2��#�;ﭿ�ޥ�܊���IA7��/D����J�%|��w�g�@^�>ﰵ��b�V�'�D����1P��I�t���w�q�AQK�ZdqT#�e�UiCCS]�(��i�]��/6pa�4[��'ry��.�]Tut��^�/ 4����G�v�y��;�X$5�[�HR�X�����؂�ױ���]�Ԗ��m�B�T����8��'���W������$�wz����e��ͅ�S�eVF.[Z������&����W��? ����h�bGw.04��2i}�/����p��@�r��p��[�|��V������[E �ob�[�0
� .�5��G-*!�$Ջ��U���r�~�3��	-��Ϲ�%��'D�B$���Pߵ��e�h����K�577�h*�"ߢ�[w�Q@_����5��+?f@���N����p�e$,�hC��%PM��+��b�՘5���r���cF�5��pa���1��c�}�.����Dl��C���}r"d��KGV�%S�h�T��h�b��B�� 	�ꍀ��6����8��c0]�~ĪԪ��j���f-;��B�\�`�o6b��}	x/�Q�4�(��������� X�{B��L��N��3OTL��!��"`����!��T%sԘ�����<۝��\��醟w�̟�b�9(-���K�_/�+\��<��g�\��4��~a�2.�6]Z0�0X�*e�� �E�Y0$��r�����C��,V�f*�~*QY�4�Ġ�W&��Ո��fL�I�&��2��y��x�s0&/6M�;u^ �HNY��ȯÇ�qCߣ\�ꎛN��)���W�Q�����?e����&a|���U.���9�Sr��i��{	×�������7�F�w�n(Q����>��/rs�f���23�3@�{���A����Ȧ{���KG&��13�\!�BS�W�����9������z
����
�4��˨�Q�g���O�o�UO՚X��6�*�`�JB�i)�aJ�ˇ��/K�ӫ�=u���Q��@i�v�	S�|�-��}j7�)8�����
9�v�f+!�����:���+��=�;� �'-�����s��8v�o�X.��ە�);29Z���ǽ�%��K�f�i�6��)A�ow 5Ƥ�Oje��
��l�L��E�d��6��N���U�f�[{�р]sR�eB��,Wb���^Y�6QJčm�k�Z�M�h�\�1����ޥ-͘x^܏|�v���,���_�m�-;�M�V�[��p��[�h����0@VZ]:��h��Wú�VNB3�|�����w;P�c�<"��� g�u���� �uS�;��h��p
����H��H��i��h�Ildҝ頭�	>�>'�R����g7���@��@�	HeO���9���������#���C���
bޙ2�-ք������A����#kN�8�����(
>����h��I1����s3�=���.�M��L4[TEc.(��t�+�66��3Z^�Q^�O�hq�uȡ���țBV}XsWl����d2��pţ羑����� 9��w �z:�8/}<0��-&.e<P�7�b�G�����Wq�(�k+:xH��E��E�4@m�$�=�|t�=6��vu�`��:q6�R�C-�!!--;o��^�v�N�����e��~m ���n��۾#,��j��ꛃ߶(�kXP��2_��}�j����*�m���+��Q:9J����>�������`�Jv���̥_6>6�����7RY,�#�'���_,T}
�xk�ǯ�o��t㙃_����#g(r�`���Y��|��U!+n�v~/��v�k��<+���S��COY���ÂP�������jiuG�A���&������^h��5
��{}��L��޳�^9�T4�儳��qN�����Dv�㘎KĠ��T����I]���b����S1��h������<�w�}�O�;-?=�4#����]��H��I��r|?L*v���[�+�}�t�=Qn�A���� yh͜(�D�����Q�����e!��V��Z�K��}l���M��'��k�xM���/m5a��U5�1�����ۻ�U�ҹb�!ϸ�И�h*�[��i�� )��L{꺴�ۊ�.4M�z�)L/5��x��fxG�r �Z���-�W�p�L��y��7�,�tt��
���-��1��m�r�,�>�F�L���hG\�>]<��~p���\�m8k�<��K�u�=�2�4sM�=J����l��ǚ����V�+�48���%�lg��!�w�C����,�l��s�*�ŵ����Lg���g?QW��:}�9P�4��ܐ)���=�����|B�dg�g[��	M��WW�>3��<ƚ�6!
��4c.1��Q?U"�m���;e�é7��5u/g	A�"�O=�#��s$=���N�)ށ��3Ieyee!�:��-'+n��V�vd�A�������	���?o��Y�;R���i��]U����&��������1�o54KV2ԉ��Euc��8I�而xq:O�I�䑾p~�C߭$���ъ�A�~������bG6a��#r]��@@����z�J�9�3�ָ�fV�Z�{xg/��@�ڢ�>g�y�#I0<|Ե��NҮH�����9������J1�JFEg ȧ�λU�tTtY-��*��+���Ʈ�����u�P��?��5d�*��ڦ�O�^ Ӛ]Lyw�b�[$x��`�3���E�J9j�2��M�	wc���_��</����61�(	���C"՛x�&��d፶�����A�6�Mx�R;�J�kb��D����xZ���ն��I���O�q��A����G+N�����މ�_����PI�ײHih�Ǉ� �Ett��ZԭN@��b�Oz����n�x{5�� �ӧ��0K���,��O�㍆�Z��$�,��h"�c�<�<�~a4]�ɣs��1Ե��4���Q��>$��x���r�N�`����I�d[�-��h���+�3Ё:߀��W:��(�yx�]ۋ]/B���_J>��||��0�L��r�֙NTZ�fqx�L�RQL�o��[̍�eYA����ew[K\��\����U����^WLe<Ū���T���c���
"�~��}�u܇1<HOZ$ʋ�����b��} ���S�Yq@�n��~AZ:�S���S�(ꐴ_�bj�Xp���EU';�C�̈́�#N�]`��Ա�`b�SKe����Y^�������~n���Sdy��hH�IL	��g���4#�����}\����4������=�@�SR���ۏONN��~�,#�{�6eBQE����G�>�D?V��/#�K���o���ד�X٨��~�v:���X������ �V���@,4R�*۳��K�xr�FY�#���p�Ȟ���q�A>�{����̾B�Q�v��C8�9����� �k�n�����s�p.*D@�a���b�T\�?�/�-Ƕ�a�����j�-43�#cI��a���/ѐ����Ċ�3��+����㧚�nb�(]� d�C4sH�1�0�$�L�o�����������`�ttt�'� �fO�� �úy��1w���yx4���������<�w���{Lv�;"Ǟ٢w�3�Tѯ!GGG�(�����q�������w��������,���1Q�`�̞����=�V�쉦��Ҳ��mԊ��#���fYF� �&�^q�P�nKJ9ҏ���b�yYBz��A��攢�XB�z��K�IE�P
�+/��x��{�\Ԛ'��X+�7�}�ǆG�lz",�z�7$�s<�6�
���E�
�=:�����y,�	�D��	�I��8�%<DP�{�.4���.=򁈥�F�v�@�K���%�����$���r����n��ZP�}8P�	�7�F9�ts�C�*��<���q2&B��[��+3dp���W�%2����e���r���Z ��%[%���,n5�*�fs��Ϳ�!�.���sԃNMYy��r���a�r�&���3=��L[�k�L�:ghp�ֈ��ce9�`I6���v�3��Xjq�e�M������W.�ܻ-�"��?*e��c�t{�	O8�������=�S~��Kzo�{�]V�Z]V�� �=�U���4����'[<oĊ����:fPj	G��	�^�\�z�4*�CB��)��uS���ŭ�����e�ڕ�r1�/;�0>�bI=8w2䲤��Ś�@aj�� k|��m�h"S��`��Y�:N����kM�1p1�b�Z�@A�F�޼OƯ�؎4��4L�*�R|\_�;��[�c��5�T��-#ٟ� ��qyV@.R-�däg�+(��N�7������hS�lo�&�&\�Ǜf��k��c�I2mL��E�`(�w[��A=�0jmp|7����u�}<��ԭ������X�t���%_�b��Zגn�\¶�
m���E�{��NL�C��wI�M��~�qH4����VMI�����b�!����?$ӟ�}��](ݯ&��~�;\�ڤ��6U�M,-`9\l��A?�I�rM`�x��Ԝ���M��g�2���� ɍb2/;��5=y��������igo?|yy9��g��\HH�aa�~�x���A�L�-괩`z�y	"xq�Q2�ޱ{�y��5�~�z���E4=|{�s��O��}���gO0�xc���Hf��,$�C�����eo��ŉ�����\'Ԑ2��e�~�V
����2`���U�/��5Yj.:1ٗ/t.t�_���~�Jg�)Y>��5yA�K��|(U�Tfl�e�p�ᷞ�S�ex=Î��GL[w%Aj�aeH��d�I/Ҭ��D�@ ��]Ɍ�qX�x���cC^�r9d�R=ɧ� ��㛘 O!�u��8���!5�o�y�N�����4|Oej�B�[]�b�J	rӵç�_qɥZ'FoW�O���\ô��R�,;dr���v-&�����=�K� �s���]}�1��;���>i�ޒ�K�)��zT��n��25�S�p��]M��u�qBC5`�F`�F?���!�
����ة=�	M����
Q-�����)ܵ�xYوp`��I���m�N�"^�)SZ�v͙f�F�ێ�A�9������pt�Y�6��#�����g�F�d���}�ݪ ��RO�p�4�b`��8�8q��>��������g�����]����7p��>�[���k*��v�~��C�_kI�˘}.��.o
o�����L9�7�۽�Q����H(��`�eK��̓I�L��u�)�J��od\p/Ur���x��ܩ����d�~e��_���:�=O�Q�E���RgI�e	�Lq�;7��P	G�%÷[��K�URJM�̰���o�k����و�=���<�P�u>֫t��هLX��`GXc�^&�>��չ����	Ҵ�ᓅ7m�ĪZ�Q��$x��4�w��$z*uko4r%�釾t�؋'Ge��nܘ���t�ޭl?������P�VU�S�L���u<Q��_@���%<�FW���47���LC�0��N��ٹ>��3��C��̐3���i��j[�T1�P-44�xKO�Y�4�kh�E�#~��:�o9��f�<mL{B|zhf)A�V=:*�r|#zņ�Z��g�j�5��>nZRɑ�ɪ����sz�m5`�`���8H�D2�){=�q��ES���S��Z�zއ!�ß���}����o�~WaЫu���|H�#PC$>lT7��^;[�7��.��Jw�����7�w{��e��io�Ee?���9e��M�.��>t�Cg]ߦy+H��Z�T��ߢ�}�O���t̈<I��j�+�$�F��Z�w"�J/�����¾4qKs]iq�^��J�j�����-�u_�
&v6B�e^p�"hG��^��f p�������,�-qQ��ۊǑ��%�(�#�x�z���()\�K��/�����XOX	�4��%b�kI����kY^q���1��te�?�|9�_s_w&�?9�)�3J̈��*K&Go�ţ�����M�-g�}�U�;���6Gr�Nw�Z������\�F�Fx�#_'7\�����=2f-?cHwf�*��jR�_������O$�l6�|x��	��ňި4�2��[=ȆT������[ʮ����`ⴒ�5:�L�Q����r�A��Z���YJ��{l�A;Y�t��^D)�9��^t# �7�͜�A��E�w�iaČ+pS���9ׇ�NӲn���D���\�L72�\pϮW��������54|���C�)�؝@oݟy!�D�����Y����bE�'���U�o7Ռ��$�yFގ:#I�f�S����e�3���}����2��ԃ}G0p�/���Ё�7>;J��	քV�Mbގ����78H�Tu.�&f����WYj�-�Z�c�&��&����ZyCȟ�{��$7i	gx`BFA�����d=za�>� {��m��v���g�����V��S�ݱR�K��c�#z�7N{psē���;���m�K���H=m�W<���YtH��ɧ��5����"��&��������������Ld����G��w��,uF���yni�,��ێ�Z����E֫8�L��v�7�SC�&f`$[�h�
M#��KK�ԦV��WeCc�:��(#��EYPh�]SC�# ���/�q:[��\�Bt���La�����-,��ඬ���@LƔ0�$-���y:g��޼nX�� �촺m?no��\J���9�X�+����fP
�!h�6~�Vhv�K_�Um��:��@q"�f�Yd��n����!n����*e�ͯv�����]���d�tW�Sk'��(8.ơ#9�6ׄ��m|t���%]r��� au�{�"���-*d��@�I���Y!�!9WV�J���],���ez�f�n22B�tI��`9������oi7��ū���l?غ~�l}�ohfQ��ѬUĚ�*K�����0�%��w'��7v��_�<�R/d<�{�kA`�5Dы|��b^>��'��e��� g����^�̙�X����-�|�3�=n�����ڤh>�5d��lX%�%k�q|���_� 94MA՞��Ӎ�FJF/���"�@�R!��^p�����w�D�eS�Yr� t^����~�Tzb�y���O�te�@����*Y���Xr!d@�V�\���� s�����y>�?�r}�e�r��es9Ye���R�Y߬���h7u��+=^�8zzH��A�u�!Z��2�,�ݲK�NM��~������U�
��j�O�
Et�i/�p�$ǔ��QE��	�|U�^���j�;�Y�ڗd^�ۗ��⚈%f����'܁Q�nEꞨ�_�D�I-�:�m��;��N��1^Z�vMp�v>.ɸ�0#�E�x�:���m��g�g���98�"�ąT���Td�Qn9k����'G&��� ��*�N�(�\Z�e_�ƽf�Kp����D���)���/ސ)eO1sH�4n�h��<���]�����:+p�0#��0�DvY��0x2��Q�aQ��Q���������r)�ת�ٸ�m����*�A��֦ȀÔ��}n�����.O�`���c�	s���$}�0g0*d%�� M�]��VDBO��� 4�0��&��8��?_E����Ă���@Mb ��K�_K��T������`3 �҈˺���H� Ɲ�t�@{�K ��7�^%�m��zBh�u2ܘE"��J+�#Ak��S��+#KXl�z��챛�3,�������7D���!�z���O�7FǠx��3��L�:���P&^AfS��ۮ7����_o�.��9"+���L@�b�O��r�9�+�/�T7Ht�J��	�M�4��� ��O��'�����?���7��|���k>7m&=�j��cS�FŌ��}I ��.�E�D|�w����FL�4���9|��%f��X%��GF�2���t�S�
�*O��g��ފkf$��3;���A��7c7G�Ub��Q���^�+<��R���N�m���A�_a�/�{͢��qn"&�;8�#.��J@W�4t=��=��3peN��(;����4H� H�?΍��_#���]��G�Կ�����^ġG%Z|��*b�NOu�0�FH�Zj�
�H`�!U���8s��X;�-��N��]��~,��e�A�>Z\��.�������k`� �Mz&|^�yuK�Z�r"���`��N��װ��h�������n��N4�m濥a�Wy�.fT4�}�K'"]��^����`�6(8�+�����t�N�h�v��D/h��n�Mm1�rN�qM����m�9u�OYy�l�AB���eT\t,tKgNzv�Fu�6�6c��<�[L���������Y#(?:}�;�];}��KߣB%D#C�*���������i~�1�k�"g��,e�/�B g�����6�w:��1����%�����tAk�?v���9J(�
c�Va�"�65�B(8.uM�����z���Ye횫L���"�v.���X��	�?�^Y\�=i���`�Ӆ�1L����+:����p��xp�z�'�y5m�sH'���C/!���)���($�dHy�D���k���xcv_�H'�j�-��Q�%i������ ���i��i�Bȁ�M���S�+%Ո2����=��c8�(��_h����Ī�%�O�^�a/����R�U'���AF�����S0���6D���A"i̟5ś^��<!b�*���!L���y�A�M6�5����6���n�#~��348�|!d?:���RD�������D�������&�WA�m}���T�X�.OCl��5돀�3��17!���q0�wg�:��L�c?w%���52�Zs���5'K�l0h�.A����2��D>Q*=�Cr1�S�_B8���ڬ��j�p|@�vy�m4�D~`퐴-f���x�1cN�A�����@�N�eQ0���o�1��fS���кj���&���O�N���@ۮΓ�F�0��?���Yj&~����n���Tr��jFr4'�M�o�`[�㩔��O4�����~�4�^"N8ƚ�c9YA��tj�;]�v8�J;V��F�c#��w:"T16:-�*"��Y��_�Z�J��
�o����Ht�d��O���FI�IxzZ����h�d�3tF)����B����QQRI�t����\Yc�� lW�I�F[4��3i����0����R��J<�}��U�$��ի죺>��e�[[3�!Д~mwU��
�z_q�!IV��-VقU���+)��Sʈ�ˑ>�{rC����n�y��MѕPd��v4���^3N햇��tm)��><�JCQM�[�Vg������K����E�z��:�������Y���c�2���aY��yKK��=W�w�l�����I�����Z��d�~��Vh'_Ot4���n��1x�!GP��?�g%�9�nBC�U;�+����s�����Bt?��y��#�2���G
�mw����ĵp�0�Lr<�k�Mx�3�\��_j'?������@�а��.#`��������
����B��g�Wv|�� ��a�Ye�'��9|��,S��
8[>�l�Bu[&��6�l����7v��B!���U��4� ��ƔE�^V�D��yf���bAOР'A��_ωe8���˦�:�����k­�`Yi"��F;����+Ү���>.�§��`����\�
 ���2�P�œ/	��x7>���4�Â�Bo3�.t�.HE�-��'''u�����VL��3�e�PȊŵ��+�T44>�Z��ڇj�:������1\-ӌp���Ə�Imslr9qJ�=Bʎz�9�� -��M����#BP��.0B�3�J*� #,,�q?`�f��>1އ��x�mꝦSc]c������Z�k���G������h����z��ޟ�Bo:�}�V�oIhϽ��i��Qz+���T�W�W}b�}ǈCDC��r�ݲ����h8���ulZ�"Y���E<�!j����_ň��!`O":���xL����v����η$Z��S��+:��������ÍvnfȂ�'8�'8ȣI~�+q*q��XF��~�ROjllo�\�]�׉!��/��ʳ���b��b��Ǟ�~a� �9�����w$qn<�><\�~v�ꦀ�ϖ��aMMML:��6͙�n��!��Ҳ7QP�s��G�A�F�D
u.��%̴_#��>��^��vv{��\���DFT���YD��EY��l�v��`�|r\p"j&Cπ��L)ʝ�e�02��w��s�m/���
w�z'v���K���u_x�ߊ��-F�.M������B���������õ�C4����hWZC��K��p��Y9�l#!Q����y�==���x�ȶ��+~����j:��>N�b��zL<���+�$�͸v�Ί3��G�s��̤2Ӟ7+D���B�h�K#˨|�]w^m=\N��>ɾM��>����;���6C�Q�z��Ř�//�]^�vޮAO������2�L!w�yTq&���P#s@s�gV������ved^|W��h��:��:�7Ɋ�u/���SC�JB��o���<��<�9�����������]�y4�����Vn�蚆�ۅ*�ۖlD���o��o�������Ғ	��`]=+��&���͓�Һl9����{S)\�U��o޼q���{*VȺI˾N{X�=K���T�˂lS�Zp�0��-@��SR�)�����N��1|	�,������ Ց���_$���Ska���\�N��ޱ���J����-������%���������������Ä"lIV\�xB���w�;��:<�lq�Yq�o���=F3�>1��C��p�i'��+~T���k�����C-_�� pn�uc�K7��u��5���-�:W֬�(���ˎj�Z���*�1v+'��z���	w22 x��)��eaƄ)U3+t�-_)�ubNu��u悫�����N;�d:���k-۽��׻�7���Ӆ
�.�������~0w��i��Ǖ<���o>�	�Q��p��@W�
����Xo)o/`�hG5W�p�~�?-��I q^�_�l��kܚ�˪z��0t����q&�h�]JK�Y�(�\n��U���m]���ˆ�u��v{��[`�=����w�7�Ү� R�� �&g�t�-+�|���5�Ļ'� =Y���N���ȇWVg��_���1��*������� ��ߝ̕��:O��x��0cx3�"�z�5��X�44��l�j�ڦ�,4��j�]};78Ҩ׻�Z]O��� �ae ���՟&�|�
J.P�"��{,�Pğ{e��f��͏+�^ZB/ヂ��4��E����e5�>��W�> ���#PP�a
I2D�H}�σ��ޢ6y��  f�'��$�
��/4�:,�^��������ٟI����l*Aw�����@���i U�-*���?f�?������RRQ���qY�Ю7Tv��y�ޞM��������N~F�cY�.�?����&��"���ˆ�Y�}W3�A��_^�Te�q�;?�Z��ФD�*�&�������E2��f_{܅�(�ō@�åG�.���X��x�uW��h����ꝅ_��������r�-kWZe	�>���R��tLƙ/{�[n�{Qz�7�R��+�+�����&Y�om�ZS��~���� Z>[�Ǧ�U��Y4���@TӁf�KE?kٺ�f/�Y�!i'��_h���Cx+gF4A}Б��3�ǜ��K|��M�������huP���W<�	ޡS��Tz��
����hM��e�:F������+d��j�j���U��t�7�~U�F�J�Az�^i�J8�\��а��[�^���6\�DRu�����1k�NO�$���zZ��ױ�d'k}7���oHӢl�����w�ݭ%L�� ��z��ˍ�K�gˑ':�&��8$z!S�qH������������~��"Y�
ۍ�3��Nz�ZYi
�9M�P6iq+��7��${���,O���8�4
ޠ��E�ƀ�J�;�=p��s'���j]�zzb����Gtj�W����k�[���A!S�\&r���C�t/baZ\�ռ��cW�ע'[��X�=��y��e7�Jx�ծ�26ڌCt�f[�� �NR� ⡼��2M�n�h�>7y5dd�1�i��֛�g`:�˗�eJى�kѯ�N_�B[C�|��l��m*Bܑ����@`2�(|��-,[�vt��;�^i<v��JD����k�1#xC�=��<�?#L�I��bp��Ʌ�m�����L��� �"����3"ʹI�4�Z������N/<��={��Z^�W�)-������S����3��ytZȼu�#ek|`aR��/GE.�L:���?4/�YF��6�.i[��q�tǻ��A�۞�e��jČ���vr�]�ߐ�6����ViEF�>��,׊���ReI�noP��"٨�;v
G/�SJT�צ�H̨߮�b)ŕ@{�.#���6s�j����K��QC�P�3F^�H���Q1��b�w6/��9�.���w�.8-�/�#�����[�'BL�5�N�ev�s(�z߼=��*V'l>E7�Mv�I���2 -�{�� ��S@N��y�g�ic�dUپU�:3A3�N�_�^,�5�L9�*�כ��	8-�H3%�!��˺f݇���kI����˜�Vn�& 4���/��.+�͔�HoR�R6��y�Y�B��Cq9t���~��������mT�U�	9��v���,f`	3Ȏf��@����s���Wy�"�h٪���9��\x)	h���&Q0cj���rb�J��Ɛ���"��~���0D�Xu��S���4h}3G|�� ��$�-kpB��[�>䥤K3(�5���֓SLU�>�'9���K<����i����o���_�~+2�{�G!�'&o6��L~�� VF��̟D���bWc�c�Kѭ8p�Fn�ܒ�ɣN쉣��੣#�>Mw�d1
�Ȕz6����RB�6�u(L@���*$P�q��>Hn;����Y�]j�U`���z�=�9������*�Qj;9�9����+��!:+���G�W�����ɑJ��gx�h`]I����C���oo6���]��q�D���E�4��=󑹽�6hL ǹ4T�M"��� �ύ´�$2/�b��� U��(��J���Vd���t:ͨG�޾7B�n\h/�_��[�n̦D"��e�׿��Z�s6����l-��2�#F����b�1*I�%���ު_��fy`n�3Y�f�	�1iZ�\��#�Op�D:��l�+5�=�n����Ql�f�f��!��h�4�e���w�3sL�0��?hܛ=�4]JTc�?R�t4 2*�_�#r��i/��y�����m}�X�k	A=�"#��j��Օ�M���a	T�Ț|5��w
8�� �8���ȗ��<�r=SoW�#G�1���Ty6m�t例�����$�E�/��n�i�XVy��M������a��!B�������U�r����m-'O t����8��uF�EUD`m�R��Wv!�#D,�r�;�ǥ�T��d{"�A� ��Ϝq�^�Y#L"�x��ja]F��7g��!�.��K֋�՘��1����|~���;��R*�a��[>MF�@�no4�9�։�ş�����WD���o � i!����-��x�Z�lv)�k��7���d#���ٕ���8���3t���s��݅� ��0��>7�'q��@W�"��K/M�mcKg켐�t浨��3���T�`��0���U���ҍ$ ��Q�u��O�{K�"a:��/��&L���R�ĭ%݈jl�.�l.f-�X|N��\�@Q��G{�b�:�Fd�3�{r �sH��'"��J�M��'i�)��wn^OH���c;�~{w��������bG[��I縥��s	{�Y����Q(
��%��dS�vx��(�������c��ȩ�� !�[v:L=��\g�0̥���sHKL|�AK:� �me�zeW�1��Ņ��ͽ>%46 �̑ڴ99��ݰGJ<D�J��Mrb�|E
(��4+T�;��[��a��I��U�C�D�F�#@�2�=��a,����*;�rG5h�����7g�#�x��s3)\~X����4������A�'���Ic`�Xn�M���#��6�}���ҟ�D�jm�X��KD6��t&���t��%UV�»A��ZE��6���uXǖ҂8��2�X�J�#>rKr��6q隝�V�MC,�X���x�xR/�g�h���9㏿�(R��έW0�˻��S`<���ՙB�	��sQS��X���.S�5j)C���6��31�Y�V�~��ˢ�z-���dt5�>b�kn�$2�<���\	�g-��@���ִ�I]ԍH�<��@���*�Ѱ���
�Iva3|B�̰�	/��b�aB�ݳ�w��2	�璒�y*:���2&+ꇂ�~\n�G�����m8��O �MϿh�Tsj�E=��Y�u-�K:­�Y1?!{V�I$��%m�#*�q�8RM�t��u��w��O�\�~X�M}�)#фO�ԕ:gq<��P�6s�)�\-DP--F>)���o��Q����\���Ä��P����2����?G(7̒ƨ���<l��)���� �T�@<��!_��;[�mO�_e��D(�`�{�D�$$��Z�˒��xo�)o$��v���c��gN0�*7��3���[		E�J���_{���} �H�Fg�����C��G(�����h�/�K��ø|�7+�l�C6"�N�8�pw�	�_S��O�w��WG|��Kh�ߐߡ��\��.���]Y(9�v5x�ܥ������O���ta?=i0TS��ʊu�7cML�AV�r)aEcwZ�9�d�+�L�w.��%��{��s���"Y��ZW�F1����������14�m�?��*(����:���Cpwwn��݂[pwww���ap��_u��i��z�vw�>���=ƀ=�v&�*�?yd�ݵU-���&��ĩ+\]SI�l���J.��cFQ{�7�k�m�L��k,�3��L�G�vW��1�7�W��uAu��0�%S�_�F�n�E�57=5�h��DF�j����Da �>Z�ξ��Yz$ӪG�הp��`0�����"ةU��3��Y~_A/G�p*��n��|��TT�^��a&�Ϻ�U�6RQr��B�wO'��G��*fG@��O��e���D;8�ٚ�M�;6��%��0�v4�3'0�ĵY�=�V�TB��DE��ʱM��C	(�������,�ǎ�(ݘ̀�+Dʨ��(�����$Z�P:F�a52�XMluB��&A�$��nݹ��5�7˗�R���Z%�~���J�o��?4✢
PUo�It^!r���t ���tk��p�=+�q*sw��ɤȀ"bJ	�yW���C�H��-
�^HZ���� �/_�J:���:����7�ĉ��Sѵ�5W�U�]��#�PAFu�y{�5r2%��Bs�E�&Q�ag6���5�ގEV��V�EV�~������ǝ���m�w`U��̕�2k�~܊�u�D1�6;ի�(��0	���t�3d�����]C���d�8�7�魒nPr��!@RK�}9�t�s��D�Q!�88G�&�Ȉ���M�(�^l���
!��U��q�h�L6�w'I?84��s[7MM5�I�}�ҁ�����z8RK�VH�,�����C�Suۊ�z���*��?���K�\t��F51�Q�^}��3X�1����Oy-�%�lH+Ww�ǿ�Й�l�OF�Q�};�慞D��T���gsV>�w}uM��(V���Z�Zv�}?���%*��k,q��2g4i3�FԳ�V}͘ݠ��i���v8���]&�Hc
,с>�0�z�����/ݏ����!tj��e#��7 A�g����ATL<-j���51Y��w�[���B:��*xB��d��F�T�@��>4�[ۛ|���z�GU��5ξ۶�⼊6`~�\QقȚ�2/��ׂƶ���ށev�$�V��~�q�o*�����7�w�_�n�;�AEh�䤳��g�?+RA7iq�/=�B�H&�4��_�6&Җ�P�)r�8%��Hx�Y5[��!n��f�l�^�H��	�/���?�~�C�U�*$�����.B;"D"���Z�*�m��$����,-*0�@ŗ���t�	��4J٢�����e�'����iw��Ʋ^�8>R�N,�QJ�L;F�k��ͽ�1��g{(��g�ࢫ][�i������Z�kQ�)���´q�,h�� &�U���l�S�vt�M��F���ac�Z[sCJR͍���5#��#[/���@�:��rN���۔�7�_�g����Q��1h��L�E�\\��əK<����l#8?���=;-W��7��4f����j�FAIE�\�D)�㧚-
���׵��/��dj��X�\����bd�N;�h��:��䃪�P�F���1)�ʢw�U�\O�j,=���ӡ_)��@:u0�np>ƈo�2RMxWŅ�Lσ����I&����o�+i�:�����F���E.���!KƓ�°F�JL @<�m^Y��F��G�0 ;y~p��)�-i 1��F �~�4š�t�Q��)�o$�W�)����#�Z���x����>�1h��^T����[�(����4���<�F��Sѱ<��ծ=t�i��xjfP��	�G,����J?3�Eh�҈�KTuY�Q/d���Pۀ�4t��w���-���>F� �%2�P$�P��#����+��uY/�	�'�����+ZI��|��}�x�.<�I�Èi����o��W������+哌�ΉՆR��=qٕv���+�Љ�4�:��� ���y!�:������0����,�k���ju�K��Q=�֠(�n)J�l�k�oy��H���8�: ���i�0�e��+�a�@)Yh�/�>��K�������ԓ�/���@�Bc8��[(@�m�A�"}�Lo>qΊ��eS���=�iLάn9}�VKc0f��jM��y��\s�������uV���&Mŀ����+�:
:�yߙd�)��F��mt�����*���ڃ��^ܱ�U��t�Q�t���X��K����}���ի��1I"0	��A�����Ԋ�?��+�k���M ����
d���d]�d��9�FG7ǚuv`���}�dp&���r%F�o�6�]��"��^m���+d���G1j��6?!S�rT /ˀj�}���ږIR��B�[wq�2(�٩ן��||v&K0XnϤ(lz'@�G�W �Bl�����9d��pQ)>'�%�?�g��?<�_��٭~���*:fz�[��Vi԰�n9��
��6Q�lj:*��w\��}ޣ���,c@j�V\ic`�q��Q����A�@���R��z��3{v�^89���!���k�]A2U�$=o�6�hW<�0ݦGႩ�)��[�̓����ZL��E�\��O��U��s_�O/�k��ᖐ�R�e��_��D�Obd����b؟���ɘb͈ަ(�����PcEO�2��
��D�;���ظ!ט�#ᘍ��i�ڭ�JQ�+�OTռy��K���ke�9[�6=!�O_m��]c�52�(�:&��5�
����@���u��q�a=D��(�H%D���>4J g�ktÎ(�y�4M˫#���"�g'r�L	������`�%��ì5�g��ڃ�#K0�����I:�8���rh��kО#�[c!P��p��&��*����~�ϞO��2؎���u��x�:�tM��#u`�_ۏ�6��!���ӽ��N:�����"]�����d�
��=�R�X��,K�S��4��,e���&g��<U�/�N�������F˷�A�Jx)�j�jL��[�=���B\��{�X�����CN? �]��F�"�����F���5BX�n�4�<x�AB�Z^�:/�?^�HD��0�m]h��J� l.O_�Q32��>ZR6��9]Iy�c��g����B֗�'�Z�H+D�{�-T��Lrp��L�r��\���M���K-��X�,��^��O�F?��cL��1X�a* ��(P:|�-�� ��
�Z`4��}�2`+{ED6���v������{�	�ޛ
:�~K֦�`(ǎ���+k�>CA��NRQ��m12�N��!~5�9�<u�E�r콸�?�Dӫ�-�n�Gwh���h�D�i��h��Ӎ�:�Z,͆���CS�>nΓ�偉���-�xj��<g�B4Y���7C�+%�.�b��a�'���2Y���'�-9������qٙ	�j�k���-�up��{&�jP��0%ǖ��)��h��9��?u�I����cD��u�'�����������|׷�\D2�����\���襪��"��潷�C>���Pd�]V>}��C5l��OE�<a�j�_3A��S�UG�(���R�}��|o%ٲ�=�iP������5/lԟXJTIfx���[��R�1�_|τ�f��%�QⶐQ��j��ᱶ���.F.�P�=�mw� ��	�&�{�ox��HIi�ي��Q�A���긶��!�dȅ���\0W�[�㉍���jO�v����P[,�����e�8(�w���J�����Sh����,Y���t��m�G��)��nC�b�����&r�h�-�Z�WdB�b3�~�Q�7�`<�^>�4�K�����c]�u�r���1F<�X�e	�z`��t�	m0�~�jN�e��?Nm%|��g`~���<�OC0+��Jj�˷��g��?b�#ihgR��F�!��;d��E1�����?��P�!� �ֱ�����q�#��W��XK^��(;O̭�>؋Q
����9�� {���x"��G����I�]�w��.�Ƀ>���>���f^&�}��K�/#�iӫϴ�!�uZJ����[%�5���m?�
����^Ճ�1S���h�CG���r�5j���l�D�e����.p���~��yQ��d�z5n���8�M��ێ��z�F�a85�nʮ0������o������ƍ_Q^��6�	��o�X��#�ok0��'/J:�a�f��a[�Ȩ�Q��'��ou4��oɼ��uK#;˒~s��f�������ĭ��8F2�A:�4�7�Ҝ��)P�g�;V���m�hx��+l�"qY]����Gm���ZLOj��q[(N���7חA3�~-z�_��j�/�Fv��s��=�0!��ٔr�ۤ������4S\���y��s������j�q&�%3�:#S�ł��m�u!W_>�l���M��ӽ��Q�2�RH���-ǀ���o���T(f�u{�]46��x���=x���c�w[i1��0�P��w��a�'��ȵ�vLh�7��;�Frc/8W1Qx)f-�-$��agb
��Q�'�����&��$y=���~s4���{��<f�D,���{c�z��k�[m)(��<p��$�q����4i�!�ܬ�	WtM��8%<�i�R$���V�R���I��������瀄�T�R,;N�p&���-A_1M��S�gp
/�	+\b�+Ld[2���|#�!_�T�l_%O,���������?�K�{�8�c1��0��� �"f�9�Ǔ��;�Gy��=D1s�d���/������m%ǆ��j�PAk�q#`���h�z7���=�3��#� ��ɡn�Wj8��A�B*�[��J��j�;}Ӏ+_��8;!4���W�Jp���4����V(���֫\��5�XhU*��qE�J:������`�y��K�X�6e�S{���Q���ڹ�|r|Ͱ�7�w+��ot�\�v�A�'�CA�Nܔb� [=ɳ#��+�z2��Y�ޛ ��o(45\��Y@ ��W -����6Š�_��7�a	j��Q8����^2b���>���7л����Ή�;��*�.a���e�E�������O��J6����7�����--�� �kv]az}u�qHTc!�#K�ɈRU���h�g�<�䲩�3�KK]�"Iʌ����^|������¤��p��H�3�w�X~�������g%`�`6�f�d�=��<�>�3H����o��#��A�M�M�T�e����o��3�̖M,ꎃ�$�N�d{���m){��d��A^�I8��~�qX�@���v��roK~�#h�e���]��|G�ϛ�j���xd�]��}������Xϣ>�2��^���	���.H���d��&��;�"36"�k����<��n-��`5��A�(�N�:����#����}]cq���3fUD�Yo�߮������<�������9�z�W�� 3l
�̧ۡ�w JXQ���D�f+����޵�K���>�Hp�
F����O��٫����(z�2ڹ��.Pm�:p�*(����C����~%Vl�z�e~��Uд��<|��e�b��	E9	���~��bV2d�?_U�TI��'��f!��{/wh���:l��/�FA	S�ֿ�?�̚P]=���h��i�uA�g��:F�epP�8�d~�����������A(F�^��$�`a����"E`j�]M!gg�������p�0�\�3Y�>�e�r6mq�FW#�Di���ol�r����]f+�'�XE��7�ig��x���L���GU�&��a�*�7:�c4⽉$�g��W�J�ѣ��m�B���*�֤��ۨy����6��v�R�$g�\�!H�����W���*��Ѫ�n��V�
���9������]	<���ɿ��yה��?6���r��9�ƻ�m�SN\���zu?w\�B�l����m���:�O���lni�ܾتU����)ﻕ��dﷁ)��!kY���,Cs"8^|�\���騙�׼S�7��I�����x���OS�H*�����&�>��T$#}ʼ�Gw�a]���T��l��w��B��і#�TD}��@Ol�7�x���b�|�u�
�u|�n��E��c碭�3W�g7�9ز��	���C��W��1���#\0��g�f�k|kw�{ܾ!ý��:�8�zB�_,�MS����p��y@F�4�m��&�M�By��p�U����s��=�U�=�QEA���q�� VO�'� {���%S;�b��h�]�~�b���#��-ڋc+#&=A�^w�n_�<k-g���@,y����`
W%;�Gػ�H��{�8�"�F_T�#Z�~�d���_i�H��Vt��f�L���\߾���Y�e�o�j��l~�XI6T@��'�Am��(		Hȝ��v�MLf�v�V$g��07�����]��&R���ﭿ��������hb���y]X�2�7��qv%�DJ�������tz(��B�`�*�l#���w&�.�M �5(�kV[���:�
����z�`�B��/txʌ즖;L"���[�f�ǋ�/��4��X	�	��t����ـ�i���f[�;���pA:*]%�Q�v_�D&�͞�)2�Z��ʣ�pa���\2E���f��ߺe�$��"�n���Ao���Ƥֿs�t��č�uK��܍��V�_�9�ɏ�{p쏘�!j��]Z	�:0[�GfǬg�3zό7�WehZ���>q	xf����ˑ����l�VKj�u��T�|b �S�b��B����ܳ���u	;|+�u���Is�q�$��I������~�n0�`���I�/��I�˕կd�lJ�"�������_��d���t8u,c�p8�7���Q��
t�Ҡ��	u�:Y����SI�VҨ���X���hn%�Z�1�%3����r������0����c��7"#
c�����g��+P^�$%7?�'���@����w��6c�I.��~D6��,_d�e ъo����4ȴa;[�i�T4����;�/����aw�y�|:�n�G�y>NUnC����{#�wd�Jh����_���� F(�)_� �������Z�1#�-�v��_֕XÜ+�躐,܉,[F�+ޢe���E�U���G�y�G���L�Ì�d�=lX�t�Y��`5���'���y�2v/i~�zu��N2��T�v6A��)HV��)fN��{�;<���V�	�M��Th��AY�Z_����o;���~\֭y�(3�_l���m�5�:r�ui��e�P=��M߽�-�g>��+��!�7��Ǣ��n���'�n�	����Z��� ��cSUoTA����0��v+��6���nɋ�E�%zX�
���ř�B��r�#S���Fc�ebh� i�㈓H�F�f��Al��L�"g����D���	�d���	Χ�7�CFA���ٚ0xc����6���d U� �<$������z_Yt��Nlt�pe��܇�RU�6q[��Fz��c���
s�/c�bz�60��M�;�(
�O� ��#�/��
�[<����G^V	����Fw����(����X1C��K�b���t�4��O��rU8-;BJ�!7�XTde�HZK�G����C{�������_�z�p��@�R�����	�fՏ��]�X�"l4b��l3���d�Q�Fj��WwsSܜ�d�;;�z腽@��a֗P���#����"�V(�~@�^�R�s+�8�N$Xp��&�� D�c7M��N�2��
E��Sh_13$6��*)Ś���Gg��H������,,$���ܯ�r��;Cf��9�H�zr��!�������N���j��FC��)!j'	h����i��M��,��{���#<�&�"���e�s:�؃9�c,?���hh�g�T�f���.����k7�-ۄ��֣R��W{X'@�����y��Q>�!�n�I�#.�!�:H�F�Ł(�iᗘ�;�eeM��]���e$Ɨ�;N�L"a4�suoУ������_������1��A#� _t�{,�V^1!��	@�`-��0�oѡd6�5��s�Oi9}+Nz�Y��H�u9�ke]t�%�H������������p��U�~5؊��l���I��8�>��o~��1��Ŝ��6b�����؏����[��IE���+�+�6m�m���e0IH���P(����:��{�'C�m!}x���"3+-o�h!'ZO�u���!���I��g�8O��~A��7@H�%W8�#E���ۣ\?
Л"u�z��Z'��=�ɓA�L	�	=ΕM�M�YCE1�"h3����y�߃��A���<���E��v�����W"��1I[0���J���#�||^	��X	���u���ͧ9����E5Q�E�U�f;1��?�e����6�=7�:�(37�+�F�l)H���;��S
�A�0������Ժ�k��5����h�^Aۿ��Q��t��;3Φ��\Q}S�*��_GL����
��2͖2�xqvy�.	��mS�ԇh'�����g�q*���s Y�f-qK2���o�����G�#����)��*6x����㈘�h'A�"Wm����W:�lN��O՝B�,m�P���\[�+�a!;8*8\M���Zݖ^��HͶ9Y�?�6vĆ�V��JL7n�v}ASR�L�~W�=Ź���G�"�>�y�r-��Yج������H1�b@���M�J��I��q+�ԑMB��A�6#�g��'���!/���Hӊ��:�o=����$�=�:����I��{����L=��x�	���SB&+�R����DL��y
��`c =V��%��^�q7�߆�4�%qj}Y	��"�U2s�y-8oT��Zւ>��~��c.���k�q�H�*O��b�r�Kgb%�7���w�]}�3\ [:�qL����A���j�|%4���S&�=�+��3Q�ݭ�.O�!_2��L1� 80�����Y����F]k�l�>H�iK]?)oֱV�(�<K��s����M1�P�}A(B�3��O?NA����)���{⃙_�)fi�ԥ�VF�H��JY�tHM�fk�#	��,�>	������]͊"��K�
�iÖ��o��A�����e,U�uY�Xm�\��������N����~/^iϥ)�&e�b��L�������|�u�i �/_��XDC�J\�c�i[U��ВDK�^wh���	����
��zȇ-/?�1CE���8=?7��(��Z�&$"��������y�J�S�c�$t�����џ?ñ�1<��Fǆb�o��S�y�pwo�(�bF;���TBa��jhb8�\��Y��;G�愻�&�Df�3���w�(SuJ�I���e[�e����]O	��yN��B\�d�x��� ��$�J&51؄)��`ؖϒv7��@h٘Ð�����ĿF��N9G��>*=�dgC�A%���D� �j��X0��)��.���.,Tk}Dp��g�m�r�d�H.���ʬ�>˹�qf:�?,((h��΃i�+K�º���q�� ����Ϗ䃮�	��}Zl	����>;l�C���~Bd��巋����a��+,�Vpu������x�?Δ�s����U�Q�& +�еY�s��[{3���Xc��4Ii����ϋR���C߫�� �"1,��ܾ�U�yv��k����Z��U�l[�G��@d@�#�ca�WDEA�aѼd)��OF���}�S�>�_���|���l7��=U�ɽ��E0+v�b!9�T�g���J�������`�F���[�1m�j�ТŬ&{��~=y�q-8#��5�p��Y8�jݾD���8��S�p�}ȇ�ɤڠ'���:�����2��|F�0���yp% �s�V�4�ZIE:����S2���`e��M���l{<���fV�2���`�F�QV�ӽ�'>��g�n�x`��e����30�6��������:> �{�!��y������g)L)U�/7�� �ߤ�~�_�`|q�x�@��M�P(�t�1 TS2��CE�`L^P^��G�@��yҩ�?ް�Ҥ�`���p���n6����$����ȹ�����ƅ�%;�rD��]�h�p?��!V��`�fK����l�:��L��4� v���
皙*�zS*��/=08%^�VC�Ǖ���V-�bA�v�Y�el�5]L������@b��
_X�%�fx)����`?����s�> 곴!u��5�>�q!&�_��t='�Jh�0��vz �+#�ڼEE�%�O�J|
����e��@�~Ș��������L�쟞$+7//���g0��*&T���*��г�]
��<<����t9��M(�������f����m���a�@(l`@�� ��a^)y��&0�{��o/u�'g�&hJh�Q	��/d$oa�?��?�|����UP�8v�ڜ"~=�w^�3<�3x3;=;3bOw�sŰ�=*}E�|S8Ĵ8Nok�g$�5$�����l�����'2���.���_��~"(rul�T�8F?��b�b�]�~>,i��5	�M�c����N����8�Rޱ�/�w����!�F~�,f�y/�O�d���=F��`џ�5R!�fٟWwU�;��=BQ���#�"�=�3,&�z�	H�[k$���
����I�S�2��S�)&�xΦ�:O�5�ݥYwe�
R�q��Z펬�5��=X �@��ѝ�Ye���%�N��F���v�|��D|��B�h@E%9�·��!��]�3�/3��S��v���I���u������	^�~�b�>�rҜ���p��w��⿐<l����N��CPK�1�=l=��o���ߺo�X��9%��ؗw?�Ú"eO�Q�`:M�!� ���?K'A|Rlٱ�
yqdd�&dy�����VvB�GL��J�����O���^Z�iDy)�R�!�
�$�ׇ�6�py�m�? ��"86:[��5�(CO��VI�����J�c�pQ��x�������=�J̵�N��>i�B Z��_��<��Q1IqO���l`<�}�*��W�j�G[��8�����e���E;[[`~ Ы���;��m���!���Me��^��Ů�ۮ��ͥ�K�;�G�����a����DF:Fiݷ�A�)}�6o��H���~��,/oO�A�O2�2���כ��Y�We�6'hXX���jް����ϓ��A;εE��LiW�BQ���� V� �($H�I�5���;a�nuu���� ���������v&XA�X�1|�k��e�)�$x���z�8t��:��#&�O���
4�H�,��U�+d~�zf�ߐ�~^V������$[��p����*�\}%E9yBbB(<T�B�e1`��QQ��u� c|��������C���Y�n'�-��fK���j�h3J�т]xgX��V�W����
͚�W���/�>`7.�v���MU̫�!O��-X���W�w��9��o�O��.1�����
r�/��@�" S��~Ԓ-�_PBW	q�6�80��Z�f�9�`�z٣��#ǲm�o��5b�����.#Jͽ�$�V����\�rZ��d��7�Dq܄��@b܅��!��X��p�.E_A�e�`<|s�s><�����S9�C
PZ�}�q�gy��
������BZy1N��e��h���:����E�_�G1��F���'�߹~���^f�Ò^4�hzL����Ӳ�D'X��/�ʕ�1�� ��3lo���"_W��
�o��vu�����؃zqC����>Bf��rݳ��]�d�d%8����Z�o/�6������S����Z�#�𵄱7&p�9�:����{p�&r�=z����|�#���4y�C��Ԅ������E���)i���w^��vI���^��txC��AZ4��&�jbi�J
cv��f��XS���EY�0�Pj*�.fq��s��b/|����&k%��מ��K��kA� Nc�!�}o�ˇnг�KS���ŧ��m�j�E����ӍF��� ��U,�&-������'���0H#@�:K"��r���� ��-V��1���B���z������ᘘ�eLo!KCX@�h�Je�E��ʕ��kY8�[5�v`mwO��������ŋ񊚭)�꭫��&$;� 4(Gew��<����yI��U���[�kn�>������[k��L�O�/�ЀG�&?���rq@�΢tÈ���A��i��L��CЭ�^{̣�=���>�K��,�}����������>)�2��,��#Bw$��NmGG���%����.��@90�������f'o	a7��!����A6�T��F�N6�x�Yku�05��_�˔�1�Cb �{j�`�����
�H�F��
�"Q|/�J��;��b~�����y���� ��@S
��E j�������[a�����1V���p��u<�S�����S1����iػ	�(�2T��?������X'5z��� W��V7�KxfVj��eh��,�E<�	�C��|�i?���q�u���+x�2��#�;���v8�]����>	� ���1�;h++��lTeI\]}a�UNB"|w�9�Ay�{��?@*6h���j=$�^/0(�����"�t�pLL�T-^@�^ni�A�@��u�)�P��`�2Z�z<Q_@�g0F�C�|(y�@�o��
���7w��b�|�����n���rC�q�Ȑ��S����#Fy�B�!�|���m��aq��}����j.�s�M�J�q[��u˦>5Wڃ���&�H�_��29}���N�3=Z�
<!��ɨ{�����0|ƿr��nS���C�84XZ4b������D�m�i5��Ā�C7K�lg�fVKΉ��e����Ŕ����PG�	\�����kb텘�g�T�ȑv����,��ʬ��B`�p��a�~��/�Q<�M�7(RD������h��PR�К�3Et?3��!>?�.m�XX�z>h�(��1F
��w��:����:!�wt��օ�9�x����x�l���LJ��	�;����A��֗P�u�ىK�2����s�,�*��jb�r�4êXs3偧����?����e���1``(�/�J�#�&���	`�|PZ�I��P����E�c��G1R�����+�	�����f��D=k�œ�*O�=\�@��@j<-RS�\bo�i�%#K�%�(�UUQ1驡D��� ǁ�_�L�6-�E��@�1�o��t)����x�!-͂y��Y��^h�+��e�+�� �:đ��rM^l������r*EZ�av��Dj_�k�X�_�;\�L ����fV��W��&�Si�`���r�DSp�V�Kֆb�R���L�i���2-p ���c<��Xe�f0�g�KD�cκ���!Vś	U�{V��n�!5~���	K�Hu<;V	�JqC����oᰘ6��&�H��d�@Xk#Z���^����v� ����7d�ӂ�0ʙq�z�����N�����_r��7��쐍��uh����b���<���Of� ��5J����ܣGLL=4�����Lx����	 ���d�'+R.X#ֱ)�Ń{!R��D�4�'\[B�q�(�u��Yr$�����>��鉮v;�R.�v}C��6>?�L�����Jwr7O��Vt���.�y�1�?�5[�k���Z?��q0fޯ�J���3���@!8��_��C��o��ߧ'�YEp�׿��h]}vѳ�9�(h�ƞ�[4k��D�A�|�e4�շm�E�Y��I��JA���_;}�M�]0��>]v&K1ч9	�U*!o���尘����q�[�����s�T�\��7���vќ�H��˵���?9��<Sn�70��4:�	']����[�,$�y-�:�4�c}�PP����\91м/otoI;���`&{`z�k��\A�.o؋i�5�^'�ah�J K	�LUc�0�Wܦ7ؔN9`]ȧE����T��[��Wi7v����Q������k�����Y"�r�]�=up.��xyp60e{;�d����HXAݿ����Z���a�g�?_jR-G��'&y9p>����l�LoBR�8���W��g�yY����2l��n:��2���U����.�-�̃2'&R��EE��fck���>t�l��`�+�Z�}+�� �!�^ݬ��X�f�e���|J��o�p�S�0\�|;�?F4�,o-����_��U���̓I.י�-4�xHH.UF�a.�[�ږ�a���#�H�%ê�N���B�b"`�����������*ES~�t�
�\>��|6�$�+k~-�߱�e�D��e��p���%`?���1z-����&p�7�M��v��{�C�-�� g����~�k��L���>ݞ� >��f�x�:ǂ w)q���c*L�����a	e�{����\���
1�2<��4�[�:]O����l�''v����'��'�j�:p3�hwܟ����C�wȌ�U]5�@8�{,�9<L(�("s �8S}o}ߚ�af�Uu�?��?�A�pPme` x󠅼��ְҒ��y�`YXx�GX}�R���J4��8�!��FA�W����4M�q��4(&'-��8q\���Zӓ���'����.xk&}�#�O���,g�of��nY菒���H�o��H| ��%���JHA8!������no!8�1�T��!hu9Rq��Jޣ`c��+X�kJ��4p
��w�����C}}��QP4��+��V���;v�J]1��1B.\����T�欙�J��M�>q�!+��mA�n����������+x�M�e����'�?(�*��ys�����A@j"�R)�sЖh�އB�Ƅ��P�&�R`Fm{�rl�RL��v"f��D^.@�f�*���EVR"@��j�����J�U��F��K<U����g���\%��i�1�9�J���a�4M����6e��-����<7E� ��������
^��� �{����N�!K/�R��΂$����5�faHŪ�t ��Y�A�Qp�|}���ɘa��A��wm>���u�t{����r����l�!�(0�Ģ4����I36<4�������I�:���=�7]+/;�T�dę����ŉjf-�)�j6e�g�O���b����eySi~��i�٦�Fv�V����N�O�\��u����'@������s{A�4����ciD��꿕����DBRJ��z@3'�x��O�Z}��1��+�ֈ@�I$_���-K�|����Htt�pJ�0���Z셴�7�1�I�J(�;b	2n�p��^�y�����(�~�^�X3�:x`n���L��.3�.�+�	�VA��X;�j�k��ĺo��vB��EG�������nV�i�]���aΆo ).��㌫x�֦���8X�+2�׺�+t��us�c���1�_���ǞR}ȝ�(--��,�����6=�eKz�VY�ppp �f�lN���m>s_,���M�U�V�z����a$�e��Q<�دJ{�J6T�Rğ�S�=���۶����$v!P�+8��K��3��S�፷���#�g�fB�q@MK���#	kl�z>�K>�A��r�>X���������S��)튐�r�*\i��dI����#�B��T>EP!��ӭ&��f%Z�y�H���W�� ^��_¹e�$\��ESpk��m���I���1`�֢����K�����Qx�'x�c���~�A˿^"�m�F���^s�al��oƀ^7@g��k�IP�Y������+�n�'��̯q
�<��,�y&2R//��e)���0�w�_��}(���Y��_����������B�;��+>;oǽ7�6�����G.�+:<�O�H�"?�y���"5��E2�W�tC�t:�1��N�~1$����?Yn
W�(�7��s�V�4i�=ؑ��B��m�n#gs�R��R�?��:+F���u���6Qѯ݋�y�1@��#:��H��It�"��ͨ�Pqu�~2����Qq���\�y��x����0��{�.����Ғ̾�OD��1��~�	��k,�O��rH7Bʂ����\k]y�.�f7�������:咦�F�H=)���z�r�k�<���4�uz-���%A�!�!��*�ß�7x2܍�!��L�A^�,���B�(&�;o��=�Z넉ȗ�)�G��ut��Hd��7��e]���?3ү�S���8?B�X�Xjꁥ�$-ܹe���V_`�]S����_Q���q�uK��ɉ�$�Q|��LtW��M������m�F��h�_8il��mL�I�6{b'M��o����`����k�u������*�����I��PJl�<��k���L3:��ъ4�U)��-���0Q[[�-D~�s9Y;��G☨���)
JVϡ'+Z*m��X�	?�q��P�c�啤�@����\*�HG(k6����B
;���`�la��`3?퇚����x�C�SmO<���_��f���{���
;I��j
�D��M>:rl��ά��=*{6I�6ͷ"b��_U�`�&��m=36�pGt�hmS��t�O*^�go:)h&s���B�����X�;^F�j+�����[��������1U����H�}�������>�$����Ĕ���8��A��&����"�^������!v���i�'0�iRL��<��Rf�b��"�%yj�
i�s�ZEk̓QDk׎��%YD�;vC]{�X��L
?�������t8I����k��{����+��0��P�_���0��֩����a[Ͽ����#�k[Z����W'ז�݉�_[R
�Y�X�~�i�P�����_j�x[�5�.����������z$:����.0BU������/SO�?tjs9J���$���
�o[��TL�L lb!W♲?b�y 	���Ȏ�iZ����h��tȨ}y]z��&j5�k$�m��xL�bԪ�2�����&�gs��z��w��c�ix�}/��
x�P�w��!�h��>�1��C'>��I�)`�����p\(���q�����y�W��y��P�:��0B�]x7O�ت��,�Ž&�����bY���r��m>��A�/�j��*���<6[3K!xK1�� ������3~�t�ϡ�b���IsO�_�/lAO��o���$$}���aذ���4�ּ2�Z	�}2�mb�QP��|ȦÂ��*&D֛lڋDƜb����� ���3}79��]��������%<ث_T5�BI������}�ߏ�^z>^HL�\]C677��)O[=h�F� �jMS�or}���ݫ�yC��������v�h�QVFl
ń@x�Ϸ���/�}}�8��AE}4&�ڊ���۪�o1Ӽ.��� t�-MI'��Mݬ��;�7n�*����1���Rm���=�y&A��q fI�P47A��v��l��a����>I�����'�����~b8����gI �dي#|���y&m�'���m�v�[�>[�6t6��^��z�`�ũ(�����X��p���^,_��;ANϫ6��5�^)���B�+��.cс�;>Ƿa��p�x�Z^���?d��4�pO��sIK���"�x5Ω�xTɂ���.+�2�Ve�>m��ԎbkO���QQ��-uĿ�����|�����:$x����+�ɴp�?��">���u5���
�����%/�����-M6&�����ȑ�5�5"E��a�����1���Y�S@_��������8;:�,W�|>��j�����3��K�_��s�/(�W�(7ҕ���+7�jT���hW[�%��#S/V�is�.�����`Lh��m��Kҷ}M%�z��J��踂#��ċѝZ�<`}�k�w^����ʔ�
��M��˄�?L�O�	`���* �τ-���o�9����ݰ�ƚ�1���8=syXu0��+�Ў��v���B8�v&#��l�ߏ�跆����R8��[�x��WH|C�ġR@�?f^�B�4�B�	͌]N|hJEU�_�d�f�u|���!#:��b �a������z�J�K�,�U��ߗ�dѧ1�]��О R��jG�c���a����u�/\���ѿ�M�^F��Ji����̤BI���<�c���mk�\��;���Jm��5��k�ѻ
���Z��P�0��r�;�ljv�������׫�V�;k��|~���杙�1�.��*Rb�Q��)J_��Ĥı&���D2K��!6� G���!q����d�W��l���{!a���9,��;�4\�!�%Y6O�bgH;�H��ۅ�ߥ֐���C-�to����o�C��qtd?�����x f����c��-��MC�����-Ú?�"�����[]q�+ö�_������WU�� �3� ��yS�b�k ��}`$��y�}��iJqh�w�G���dP�P;�7/ ;���R��@s��jW ��:\��5�艘����>8eG!�^�K#5$��ҠK��X�L�	|���X$$�[k��ޘ�~�>u�oO��^�sk��\U�Mk3�}���Бv 4�y^y�{�#gW��@g�o��+���~]�ӊ�+�C7ާ������뾂~�p�⣠\Y]t�&�3�2.ڝu���c��s��dc@������o�����z�K��뀔pR� >��? XpP�b�T���h��N�]A�B� Ka���Q�������6���O�������J[{�;}�G��>AO��8�W��܄C̺A���#K�+a_�̓�3L�C
�t`���mI|��^1��$0��E�b�F$�Sj`:D
7�h�#x� ��?�%���e�>��XxK�(@KQx�%b8��
Av;5���9*����]��-0F#h�HR�L���RR),���O�_�T�;���QmN�����R��L<�����]���et�stC��!�/.
裌q�����f�5@�'�Pc��m�R,ʍ2&c>1�\��P���խU�z�"�MuQ9�����,��U��l���G6!��%BH�]��s2BH�XТ0���дC��ޯ]�՗���"*����#Gp��/����Q��@ ��"6nY9#<'n�,/�b�s��>A'A���'��P[���/�!衾�������YФ�v!3ͥ��R3G�:3�f� YbalRRe�\ȱo������kY�)��f��H�Ț'Ɗa� ��|W��-�x C�����ڙ���Q�����h�RFF�Boo�f��#ɷ"��[4��0�7���)��q>_��H�~�i����5Y܍T�7�5SbvHp\��L��HI�r���_��2�))P`H ��b��#����:�ۤ�9Җ��VY�ƥ]�[�*?r����ƻ�|�:R�H0]֬��X/�dJmSS�H�/Z���׈�\O<g�GkԤ��_��1����]��H'�C;��G��`���F�2&��G��T#��$Cw��&]����(!9p�o����Փ�1|�`*�o��/�j������'��,X�x����C
ݤ{U��HvF�6���$�U����=ZY_h
��-��5�@�Xb����4�L�U�]�J��8:s��J�V7�8�	�v���+<�+Z�e	�0��}��d�~3��%�L)VP-%�'�	���^�*@:��Lѐ����R���-ŗq+ׂ���}xa��$[�����M�vO2�='��z7�8��닪',H���P7PW��}�	m�w��n�I#?�	
���m-H�"�"���~T��E-���� 2MB�d���0@��� î����Ǘ;�j�G6�Rn4%a0�X�<��.��4�v�&�~��Yqo��e�6LKɪ-�ͷ�,�H���
�cbQ���K[\3����p<x��a���$lf�/��j���.��Ț朽 US���)�v�#�8�fn.����Q�_�d�e<�iT!���NM"��C#	�'���A��0R�W�!���8���k��̍�SF�����F���{a.�}�����F�����A57���*��؝�_�c6� ����.ܿ�	MA_����u�ign:��{b|���:e��/qn%�{zbqv��9I�p�?A �|�欙#7����Y�zf}z{�J'J��oGŚ�>m�TI��Ǒ�]�V޻�����I����hY|ׇ���2~'���>�r�E?�Z`�=	s�{��� vGR�K2�����f �'{�29y�K�19�,�JHc��%k���"�҂�~�đӭھ�"���ߟ�:jr�G�mD��!����f�J	���""���60��2S��0y.�$�#��?�.��҈'$=�\��mQ�;RP9�*G����h'�h��-"AY�r}�Q��&�U��ɿ�l^�9��Nm-'��i	�D,Ƭ��xr$H{��F롗u1�2��^�3��j�'�q5�Q]|�o�I"�@���ˎ���	e"�~!�+D����}�����ב"�V���}W0 [V���:< J���x��ν1�~ �J�*&+@�h�mP�T�Ȅ���~Q�G]�p�p����x���}�7�&�q*2�0���{~@��צabj�����&�)
�x�W��ڞ��)�؟j^P7����xu�T�h�<Eè8p�4�#~ո������s���	�������*ڄ���Ql��МS&�,�Ȍ�_�o�YNT����)�J�d>Pp ���7��b����!���>H��ec����+I�^hL�=x\�"7�+EJX��t��u�㮱@x��a8�B+T�]/D���~���2"H��:9m#ʜ��w`�^BB �22c����恀������f��h�FZ��4�6�Q�׎7�lz;��{�Jb�IA�uֹ�+�������O�t�Y��wa�ïa�Z��e*�(Ǌ�)V���_�2�O`A��|8�N�!��P1
Sm��Wb@4Ǣw3jM	r���N��|l���}�;4�0F"�k�m}GFZ�J:W�De�[��UKhA8�WRA�"� �{a̰����L��h�!`�e��:�cg�<3>�s`KAhfgm�%P'AFJ��
R�b%�Q44^�;���:Zx�"�3�dS��n�UG��N�E��I@��A19��O���\_ގ6���4�"e�^�D�ֻU9���m}7z�/x��1/�lmNbKµ҉8��'�%��R7�����a���L�7g+<k��6�}��_ g�C�������V��[�)@�*�����@���g�aX2Ub��˺�������wj��&E�7��^s�L��#X�B"AÖ`���bZ�A�h�~�L^bD�􂈎S�+Gz�m�ֈ1b�l�)��<l�>.y��~��>m)�Q��IND���/-�N*�Q���o��o�������� @ր�Y98"*�����T]�զ{W�`ٓ����WŇ[WM�kbg�~��&d�ϑ8�*��ߏo�h$�j5��+��� �"� �R�a1��`2��\c1D��j8��qX�h��;b�_���rļ���g�N��kA.�
eqש���{�� �R��,��r*��,���.�vF7�ʱ�-�b�GB��)qD�,�V�yJ�(.��Nű���&ݴ�w}��A{�z�(5�ڌ�@�}����\*�ؗ�t�9�.�c`<+gj����LK�>Jo�w�-YG���!XB�aX����M4�0G�1(�Z�!g�3�QN�e����F���<��%�c4�Λ�bF2��khn�C�6Z��@��\М�]��C;^TљՃQ/��D�@�����ʰ�>~���.��4F2f6.Á��y���q����;M<�
E"��ǕT�����$��!bBK1EuHaT=9��ƕ����Ik�cx��z�.�	�LUW1։ ����]P��5fp���^dW	"g^U�y�3�|��]����]��� P=jz3D|�j���/�ZI�+�(@���/w�������h)�>���1%fuFxY�V��Ә�a�L�eA�X����D��1��X@[��,�1[{[1��ԇe��,]��,d�a��<D0�v)=�m���k����+N��2:V\��tM�N%�c��
e�q�a'�|�ŗ�򮀚h�q�B��A��j�փ������}>8�J�����EZvڜ�C��5����21�X8��W�&�I�+*db�޺�C�M?h�S�"�,/��R���ګ�<+��;]��hԑ��E�e���9�~5?- ��w��Ӫ�^s~���ȍ�S�x|j�cG�t�u�!��z��J�~��"��������K�t	�Z.AC�%��߷�A������cu�v<�7�a���L�r�$A4�ᕢ�G�n�["c����.�.�D8�Y��ߊ���,�N-M�:�ؘ�,4�E���I\�f��F@�Äco�Fb�ʧ��ql;@a ��:WN�����2S#���=��'b��J-��hb����7�sS�2$

����|�/9�Fڦ��Խm@�߯$�O�Aʍ�?�X�G�};��[�=�c�1�_��0��}�|�E�u�N�8D?тcϪ �7����5���/&�8f1�Ɠ����Ͼ5����>�m3Ek��h�t��ǐ���LNs��rŵ~(,ӑ�Q�0�q�0��ni G�*�efM[�[�}�P�1B_�ҿ8f@?.
!j!K��Mg�,Y���8��7���9'M�[6�ǀK�a�^vkK�Obt���p�2�a���(�~}��t�R���Փ��ұF�q��x���[��'㭾���yj��Ah~Zr�O@�f�Z�u����.�Y��a��k�x��I��R�K?�q��@5�ClKI�I�jҪ�'�-Bc��k4��Bxs��Bs+��0M=L��5���������8;�k��Y�g�\�lr��غh���X��/�B�����,D�$Ps�
���p���l�rqgT#h��'v!>���tm溚�<���� �'h�CO{�u	���AH�RB}��8��b���5H�r�ؒ�$1����b\C�	S��k�2��V�}�����s�u����t��ױ���9}�!@�u�Bѻ74_�\[���<����ټ�}�y�|�,�^��('��ʢM,��P�\_@'�-6�c1՝����0B��X�����(�w�u�4M�_���ǰ�Ú��9��Av�k_����⹬봆+�<��0F6I��Ga�����P��IU����/�6�<M��eɿ;Y����tY�=�{�D�0�͆��W�W��V9m������Y��X?C_�c����l9bѻb��T�pk�$�Ƞ�(V}�KuC6n�3B�r��n��S\ ���h�<�c��̜�#A��t�PX�|��E�n�G��	��͘<�#���GmC�� ��8��Ǥ�iO�mr��	��`Ç[������1���L���̸~��1��J���K�$H��}�ի'��2f�����a�E�p�M鑛C�6���3^&��*��Z�Jh�6�a��1��[l��;�z�vkM�\��� UQ�����u�J�h\$z2w�ā;}��ww���U�;?�r9�v�ҳ���_���SE��-����{wD�|����?��J��P������e$��-T��1K��B�Ⴤ/D�[n%���/2�ؑ8l%�t��л�L�������5\��D)ڹB3S?<�M#%(V��T,��Eȭ���B�d�߼�&A��P_Y_�;+p� ���;'�E����9L�l/gI!!��ۛ�L�`�Eu�Y�<�J-;��s��� ���N��Z��z^���d��P&�*�9yp���T&�"�7	�L;���iZ��R,o��UV[�k���d��	�z�n���z
���{�v��=c9'����<c�{�>u!rC%���0i����F
����h�&S�i�Xu�d*���e�0��Nvßu����R[�au�L/�:���?Q��a�����@.��9�G����27Î�4	�߹�/�Y�������Ǎm���/����e��6��������bl�&ˎ�9fވ��bP��u��F�$���������#z@;*���o)F#�]������?��?�.�Q�fu��;]{u�Y��)�ƍl󥒝X�8��z��+����a^����!8����7OV:�r��A%����Ǽ .͇����N�n��-�׋(�Sa�� ���q�#��<x��n='ڮ��N��1����@��1�)MM��+_��-L�Y����3a�1|(l��S���׳阋@-/Y/��Ɗ�~�0��'�ԓ���`��G���_������%��Mw����:R����ǯ'B⋩%3��) "#����:GoU�_y��㣸�OHTƂ�۴�.S����|�!�~=~.���q�_?C�$�$�[��n�r��.)����g��\��g^
f��]��#����[��8�GU8P�Q�۵�M.�61U�/�azcM>��w�~s�z�$��E�>h���F���D̆yF49K��܆c΢R��R"�0�3w�Uc�3tX�u���&���T�|N��7�l�2����#驰�X��$U��sW �\��3�g��YY�v*���;��&��p�j�3A�;�z-�.�N��$�h���=���!�����kIRQ�ѣ��@x4���ג1{{f�4�ct�[�,|�[�E�ñD���3KI�K�a���)z��c�SހW�����`ə0�L��O��_���ܥ�a׺���l
B9_����C,��N���V��g�~����b��E���_�q#Q��Y�;�Y���V��i)�S���,�B���**�~�Gu:������g�r���3\�����4�^;��g���|��.��</�^���L��E�x#K���Dl��>�~}�D�9�1t=�h_'�0��gv�)��
����_t���N��)C'$���W,~��ә� IHw�T'#;2s�:�^����sԽN�a�d��*���m�豐��}��I����J��a�y44
z�k+���n˄��ve(�A|��r	i"}я]ѷ[���ݣW��?k�v*a���ñf ���̪�����ؤ/H��v�v�X	$������s�i� .G"�hB�
�{�R���u�����P���9D�Iر4���Z'�.EwՌ�!ĥ�r��;�3�����L�:��]>�i��u��F`c����g��*F��~o��h�A߭�9�]#2$�Q?�3:���������u8�F!S�F���&��6�y�$�����>���Y�T�6�$���V��?{7�=�Ȏ㍑����oF+tkIp�=�ܗ:d*NDSb����D���*OÃF&�V\�R4EOMJ��<�{Bg9��}U�^�'����*i#�q�}���χ�kMs{v'z���[i�]�Ol��n�ؠ����Y�������~ܞ��Bp3��y�H[�V��1���;N�7��� NS9҉�7�,���t�`�`�h4�N�öB`�4�ĳ7Frj��0�x�[$��ڮJ(��oc��t����
M۪S1�/���DS�N����3�R[c#
ʋ<N��2�"�Lo]�\�a�+*�r�4�uD�F1��W����ف��1p4v
C���Q2h `����l۴��,)���C����Ì��5�l���)Ѐ��:yի��oO�:�j�أI�|p�]#���5�k�k�o���e�tA�!�\�!�>O��+��܎��eș{���J�G��w��G�P����B�'�ieЛ--،��+Q�J�Lu�����@�1���n�ӫl�#{^�aD�����K��q�sv��wx8��Tj���(��._�5�T��b[NT�πE_�֚/�A�uF5/31̤+vM���n����ѲKG��N������膆��ʃV�����KK�i
QKi_ݼ�Zb���/8��`a�rղ��S|�~z�+��m��]�ُ��&�K�O�����EEfR�	j�w��m�+@ T��=g�Ri�صX���cf津�g��[�IB��������y�GVb#+l�]h~�W�4�8�
��p\�k������I�L���I�/�f"A�]�ȉ���ſ�e就ݜ�A�#CÅ�ጿ��?S�n_̈́2M�����D��H��u�d���B�2��!�����m�֠G������y��z�HLv3��P~F�!�A��G_�����[�G��#ه����fm���;���5��vyeV��Q��+��V2&}&��蹢���b4�D�7�:gSM9��$�*I����lQ�d�^��H���r��r�!d�����$B7��f`ϋ�G���׏��2߷�en%�q�Ώ���V����g�Ը�e�a���c.��^����9N�օ?�ut17)ǜFˆͣ>_���=ʲ��w����u�:�h�"mc��Qe�?I���Kx%X�Pvks� z�������Ba{�Oe;��X����+&��2*�vD������]pI�hCC9:e��%������x��D�n8�_z;�ms�KE2ajM4������v� ��i�
Ӏ�؆�kP�̥-���7<u�>��t������mw�����aW��ɨ5�*���:ij��.O޳��N��?�`̢�1��]
0㎉��{Ȕn�!��֑�Ë����"�d�\H���F��l���#���cx=Da��;D�f6cK��wP��_�����<�EOϞ����U!�A�i�f�#�aN㤵��
BSL�X�n1�z���P�g�	)f
�-�#3$l���e\���c�lN_"�����T��F͟@����)=�t��{�{st���,,����%e b%���֟6� �\��&�K�3�G�@4{�9p��evq���5p	��v�DT1g��v

�5)�,�`�}vN�����oC|�����O�i�4J"U�+�)����у��lp)�s+��H�شe�)3ѧ~�|��(%h�:��C��9�-I1�Z��5�":�* W�����;.��hd���V� �)\�b������PTYM�S`Cu��7�����fK�o�U��W[e�?��`*�e�PҙqI�����3�F$�*�,��X��?����oo"��Z*��?u�Id�8��J	�(p�	�����~�X#%*Ճ�k��ڰLh6	C�b|+S�uꥩ4k/,IYZ��Ȋ���gpR�yb1?o�^ i���1����m�ZÔ1� uD;�E�������n,���ď��$cD��)�
���A�u^�i��ғPDH	�o1�m�S�p�&����sլ�sT�&��4O�Y��U���P���nZ>��ɱ����P(�*p�������"���W���u�����yE�l�aX4{�É�fA�ia#q����/ͥ�$]Ȁh?I������;��]��d+`���ۗ�������?�#Ucڈ��X��!�&��9i\^�b�Ht/��O���%�v�Ǵ a�?a�ێ���J;/.�8�7�.0�`$ȳs`"��7�fR(+H��W���M�5�������G���/A�r�P{{�0A��C�����3���Q��W���#i�M&K���id��5���Ɠ9�*��D��V���h`�Eˀo�LFZ��Ob���#z\VG��*})��q^�5g���G�n��C���� �SBv0�I����վ��x�=����8&�}�=2���|�?�F�3�C�0^^8%�����m5��EF���z_@[�(V��D����v3hx�b�#m���S�5��4�u���i��L �6���zu�Zh۠ �l���uI��K�Z����1����>LI~/婩I��bM ��-9.%}{~b�H9��׋I!j��7&�y,B9ݾ?Ĩl�d�b�R�H�m�s���/̲e�aG
Q7:�5�����<�]�]���ֱ�J�{ٓJ�� �3�/m�kU��zt8��aճ���;%j0�-���r�D����HM]a1mi�=�-�',<�ii��H1B{k�.'�;E�$����a�-�[�|
���w�r�W�_p��t�JI����r۰L�b��Q�����<��V��n{&�k�PE�V�����3o�\$��˅�mcP,����T�4S�؀��
QpUSb?���2�9��__ކ�zA����qu�_��(�W2H�5�X�����!�Q]摙��KaƓ��v�޶Y���K��J�P�M��PF+S����t)zϮ���8qT������@��A�[lVÿ�r�n�y��U/k	������WRx�w���}[�m�WVQqB�Ӫ|������+�|(��\	7/DW�>8���-ĖL����<�R�z���,,�����)���D��#0@sMl�ي!આl�Y!���Sy*�f`�"y�cg1.�_Xe�����p�����+ٺ�(Ea�x���4�2�u���~�ƞ}f�rF���4lPթ���͵�Ս��-��l]IS*'f.h��UV>�e8D�4N�U&�zK��7�n�r�]4Z��|#�Ҁ��8]��ǭ�L�7-�����%
��'����tya��8�S!�Sc��;����fNfQ�oW�Z�N�x(Ipz�^>��[/;���3W'�l������?�Xj% *�;����敝��-�y��~��i�&��L;6w;-�t�E��a�fmq���@�R)�T��9���Z��C��˥������˅{����B�ڢ[Oϴ��������|WLt�Y�(�,��Ѵs��
}��[{����{`6/ED�di),�7��j�g�nq��OMCh����뽑Ov������؈�� 44�ts����?Tk�ڑT�ջy�9 ��1��(Є�s���TRRG��`�&3pf� <|�c���;�_��yRg֚aq!�:U���Y���5Ռq�x��g<6�l;vr�<��Vu��,?~��w���{���kP܆��l�ļN��9��]v=�^n����>ݖ�ݢ���Azղe�8^W�rO�B�47�����}�'��auA�"7�]v�Z3�ɿv�����Q��jh�,����.��+Z^=���äNg[:��nՖ���?��c����:�營V%����5�����~w�G�vC�<�ͽ����gɣ���!j�>@ҭ�Mi��7�r�^ۮT�$|h�+�FcW�⃃|1wT73��d݄�����Ҡ.��gFO���)��BF�ǻ�)v��}�R1@b���xۻ<t�
���*��}�f��Uzv�}���ߡ��I�0���A�O�����c��[O�B�����/1��S���<A�˂�RTb&�p�\�:�C����Q��@��y�����/P!j���e���-/���>��E��ʱf� CQ>��b�q����%�DK�%�Td�̡{\���#�>/��"�Y8ڶ��4k��H^�d��e�(gV ����Iߐ���p'�;�f8�1��9lR��T¥c�\]~:�c�-,� 3��'D�|hƻЍ�T"%?�l�SL���r篈"ɭ]H�
�N]B����NP�,A��g��O�7�]�yTH��^��B*l7�b)��x��&�Q#ZƓ���҉�Y�ʔ]��j�6�D���n�נ2xDg8ػ��9�
�E=�{b�@k&K�F���ttH��4Ҧ��Ю)ϖbsc�d���@���Cc��]�@�j4�:0w�Pp_e�fHP��58��ղ��}��Y��_�yt�F�ׅ�Yl:�#��Z����G1�~�lr�یQ�2kqXy�;�k�<�ռY�
�΂�h�jmj���@Z6i*_���(�w�@�$���gNWPVV�aM��X!��'�1��UP)o��=35׾+a��3.seV�UP"�v��YM�K��B-T��L�ƦIoG�\B�so?��c��%���p|9�x���Υ���ܪ!#�%����R4�������������/΂	�{[tYo k�ѹf���F!wD�fO	M�뭧@C�7/��#C�����ݲ���G��z����:WF`��6�iw�.q��v�rd9�����zd��^*����W��؄JSr��t�r��� S��8��j�A���"͜O@�Vf��m�D��"ҕE�/�%a��k.�L��F�?<=3��P���:8Xכּ�TR�QgT�jk��U�("}nZ��r񌬪U	;a����lc�ݛ����]����?]�섓9�:Kl�jP�S?�62�	��v]]�ON<N���oF~r��t��F�K���D6� Z�ƪx�V@@`�:~�b�=Z�žA�U@PT�Tz�G]�o��W�uzp���n�̕��LBU##L�W�d��7ED#Ԙ�>�����Ŵ9�^G!���̫�K�h=m3��1�(J�U3�U�,E82���@C���Ӽ����:V�<;~C��!��gz��)6y;9�\9]�4��uan]�5D���Cm�.p�)}��	�*!
E��2����FS���������,�|�2��?��`��R����}& ö���\�����<GC>|ܘY�{AwdM��d�f�/�'�G�T��ɿ6�����?�p`�^o&�@L�T�n���[��[bȺi�c���|x{��WdK�_m-qU�%������PX��7�hs���ܤib���wֺ��NFin�VM�<�X��5���/7�s�tBڍP	�bщ�HZ�^p',�fc���-���\����h$%q��%�ÄJA!S�I#�d�lL�L�}|d`�n�����>��U��]�69Ca�^j�GW�wW�׃���Эv��J5�w��Q�Ч8�zX����6[��l4��S׆F�X��:�ᘳ ���Ģ:&q����wb�$��S��F���'E�s��EĈ����u>Y%sM�Һ����?lZ
Z2#R
���<������u��}9�;� �L�F���A^!ie$R�Zj�?�?��=��RB�s�f��*l��OԱ�S����qeM�ڝ�xw�۴P��i\�b��c��OE�}����"��,�I�H�0-DB8���:�#<�D=��7Qd���+��ܸm�� ��A��)�{�s�ە{y-nu+�����v̖���\No}���������g���0��Fu^b8�Y��u;�.�ы��CT�6^Y�pZ�7`5�e�˥�+��M �J�Grs���X�T t�.�X�8��W�i��ъ=�麳���{�I��*�[��c��M���y����X�܅��bb�	�5��Dc"�i�O��6�
�(����b�Fx��(�tmH��d��p��d�u=e�;�ݳ�nՖ0m���d����/��x��g���]9u�oII�8`|�Z�%�m���%'ɩzND8sz�2'�2�ԝ'qӽ�s0�3J�� ���B"4b�j��3vG�g�n+����'�+]ҼX���D�S�t;R��y���c<�����N�ۓ?mՇ�>(4
v�q;�3}�+��N�)6�5�R����T1�d��>�6�����ޥ+�6�㘚�pQ�ı�,��ɼ{�X�{.n�bA����ʪ�c�q�˶3�+ø������.�B4nY��j>��mb;"���|.#i��g�z�:���m��y�y���cy�P�۵�˺J�����r%^�,|S]iF�j��Q�F���C�8Ia����ZK	g�-&6J�ڙ�7���D�,:���W�G2?(;�]<͛l �'A><�z���[�=�J�%V^%u捬4:	��~nUm���Ɵq�Ԓ�!�ߦ�"r���dm��9'�l2�S/����d���g��yZ�|�2 I	M�FQ�K!��/+W�A^���u�Y�i��I(q��.�j9H����]��Ǆ��*ɇ}� A$��c�̆��5-Ӥ���QƃNF�Ep*���\/�)U޵}5�����V.;l�]��:RKp$�q	���R��*�����V�Ͷ�� ���tr��$.��F��Y-p�ٽy��Dt�Jʎ�%C��_w�s=.=��8��l�.�\��k}���!YW��i1���Ԏ���\�7�1= �PX�b �s&��H�k����Y�sc�13N(&��Ϣ�J��F�I������Ũ�������NXr2֧�(PRx],4~�e�_o�MG���¡D��mr	=M�quMɞ� �?�����p���Ĵ�6��p�vs�����5���:�����8�Sd�Cyi�1�5���oP�1��Az�=q��h=d���s]����_A����!m`8�Ik}{W8�TЭ�{W����TE,��Q %�Ӿ��BU��/v�t�Uf�=(�b�� Z�?r�}��(�.���������/�]������ ��T��9��cks��7xw���e���"�q�]ڙž�kzh�XLp�ia�\v�'�̅�������_
���fKU+���utv&{�
���&�*��O��Y���qď�-*��(��M5SV�/��_�Tm񐀄������S6~�������?�L�d��Ϻ'}V�9p'����j�d�֦� %V�k�㭭`� 6��]bMy8j�s���UqZ�d$��0�<�Zɩ��;������\E��&Yê������`�a������K_�W�5���Cpww����]��;�a � ����W��]��z��#�+J��	���<c�ѵ0�y��t���_���x;O��![��ö�@L�q����«��Fî��{�y�5��7�6a���,:�0�ӯ<�ӫFJMlte��űFY���q8�5�5����)*�R	NE�Xd͝&�C��ʂ��!�h����h\���Xu,YN�L�'f_}��:+t����:l��	��N�%%-���F�	�|�x�����e܃�v��5�9�G��\����m���u�sd~�>֎�dgj׋�s��-q��z,��Ֆ�?��M͗f��:�ˣ�%%Xֶ�;=4���)��6-�:���P����L�6�%(����r�f��f}g��9�l�U�F�=e��SU�1S��(�t�ok�4�#�Q�=�M����(�!�TR{V�q<�a_���ְ��~�V��5��X]���B[��%�m��5��h����D���$46���f������4�k�1�-?Ut	���)���:�u���9�����h�K5�ux��.b�X�[�I�4��$�	�� ���;��x�o�C8�M��ɼ�+�!N@*5^I����c� �P��"��6��z27�4n�8��@����d��!��?�o��Z�N9�φo�ʀ�ݮ�����{�>���o������pUYTB�	598s��/o�|��#QITc�P�/@�
 �oر���(�P@�#��Od���:��1�/��{�V�]�5���V���^����'�B<;�XY䉥��RMĬ�o��]�ޤ:�>����,��PRz%��!�c2�܌�VJpt9�K��ʡ(ߵ����no����84����Y���L��Q��*)�d��$��L�P�~��|�5|�i{x�6r�zz�á���帷f�m pnn�y���/q(��W�I%�U�����*/�sm�U�]������c�l�����4,H+��^�~��W'\ds���pzB���9�o�U����~L�6�ڴ�\T-s��}/!�B�І~�t�D�~[o��2��
����9����[�WaX�~~�3�ڜ��A��e����&&��Yf�Qe�®��*oJ>�%��N�&�Y�-q:α�){������Fr䔿���٣|�=S\���gt�pӴ˞��w���̉��k��k+�J6g�LD$j��O�D�]/u��g;Y�R�y���x{M����5hS��JI�5��S�e@��*�K�YĢ��pv�Cߊ�k�]u2�PX�����7]��������7i�6��N�[.I����p���{Z�)f�da5��t��v���^O��ėm�2��#(rs{�T�4
g��+��]�}��ag<��w9��B�'��q�I��h��ƒ����Z��ʱw`�b���E+�i�a���;]qX2F�q� �vm\�A�	�GfG�����%��o=�wz��Fܣ��gx��A�w���Ra�rw_p��E�go����_f��>]�.2EeʸE4\n��
���gp������ɹ�Ţ8W'CB�䷃�q�i�u��2�1��j8w��6&i5OtU�M��׳���df����i�<t�4�a�{��v�ӎ���a@� J�xަ�A��\�O ʹ��G��I�eAf�.�a%~ϐy��n�p�N%S>��Oqx���� ����/g�ױ�/T�oS`ɪm��a��x���:�z�۽�jܥl��!�UC����_��u*�[y�Tݠ21���6�4��uC��<>.�=��иN"�1��[Dn�ִǠ�oҭo��3����|�d��73Oh��u�����lN�������IӪ2kP���K�̐�_�����^��y���è�4�QȲ�fh?��Tc|QϮ/��6�#�����$�%)�~WS�W��_;�����?��F�p��
�n�rY�|�%�՜��I�{D�8�rZD���i���l���l���*qcoV�_<��#1��*
ɲ�tB����{�L�!ʪbŜg��~�K2[r�<,-X+%��}lyC������(��VB����x�J��lZ���
j0���J��PPq�$��JǞ�u�#���B�m]f�� ���e�'�X[t��2����Q�w-6V�gx������wE�B�7����؃-��F�6����5���y؜�i�m���}c]m���ֺ�y|Kg!m��~u����K�u�����[�����V6�/�!9)�xC����딪c	����|�5|ϕ�����ǩ��]�����[7ĉ׻f�n8,�5��ر�긣�s�#x�	�:�3�_IX9�T�E�lcо�LK�>��ٲ�q��, K2�Su����[����w���]Mb8Eu7�]�C�0ov�
�{�˥� e5
����Cg���b��������49����X'�(:���"���&������	�����l+�����H�#��Sh���a��-�����t\/{
[��G�Q�yu��K�q�W��b�d���[�`7��>-@�,��H�����k��r�V�w�[�69"�K���Jc��׭�Y��yi���H�[���(g�^���&"��k��5[��طN�D��Ξ�x��,=!���O \����U'+��Fh�[�R�4i,D��_sp������P����tL�4 2����=���]�܆]:`*����k�w�C#��Vp�{����'��������N��AB�ʨ�U��P�-q4�}�T �*ɣy�w���c�����[y;��ۈ��J�
[��r�(���m�V��f��2��_.Ap�e���.&�G�ߣg�^)��#�'鰜3e���x��ܻx���6�=�O�Տ#�I��g��O�Χ�/�??=�D��a���9Vt�R�H�@��#��?�'"�e� �{_ϐ�8�#B�6�M�l����+�D G�jS��調�-D�����@��g9������n�CVw���Eg$��i�����;�<ÏH݉_�ֱ����!dzF#�b�~:�Ҽ��x@(|D�{�!���\�?��{�g���	�m{>��=��+��J֧��z_�~�AN�����
׍Ⲻ3`ko�--$~�5a�t0���\׀9�twM��� �i�"8�p��J��<'~�$��H���Ó6�a���ԫ\&�B�����h�21?K~�g!aE�X�I�c^S����esǿ� ��ֵ�����#lŰ���,�
m�~���tD/�����q��X��`#z�_�bb�&UL��e�iXP����/:�x�H{
[9��jnR����S�6�۟���q��s]�I���rc����{�kv��G����:�G(e\{�,@�xfe�\��t�.b6r�t~eYµ8�P6vt8܉���x|saL�2��0ɸD�oFI�z�bX����R�����W��w��[f`���]n�	oI�N�=eN�h�,nբ�;a'0�r�g�5i,��%��i[Q���OR]5�͋~��W5�*Y>�����mȚ'1�|����^�}�.[�k�WF~��&�B)Y��,zl��Tr{����:Y�;���:ۘ�9^���9�Jؔ�Nn.��~W\�9W��S�����mhհ�	V�b/��;Db�9��-�w��~��8����: �i�-GJ���i��A�ܞ47�	��!vz���K���m��Hgw�����o��ؙ�΋-�y=�����1|���H2X�h�ߝ��{�E�ki����Ջ�پ��Z�:�>E��n���H�(�ff�9?��uZ���8ű����R�oE��X���P�g���5��c�2*����z�C��c�]�a�)y�˼��������c�k�ux�,��IH޾�QCR��/���6,��oKch�tv��d����t��?6o��"��K����te���4V�.�B�N��K^���Q%na��_��Ӑ����l����Q����x���:�G��E�w����<q��I3�Τ=;WW�>L5��zL�iu2���_��0�9�r�59��d࣮��_6 ��}��}�~RrѩH�Oı���;e�ɞ{G ͎���6�L�9Bڙ�H����<��+/�8�RkM����ߩ%7���\��8�J$����t��b�����me괖za�On_1
 _�n< I�����|��B;M������F��׉��V<�p�U��j�0E�����gaJ���8Y:ίH�_�K�SS��S���zGA<��t:��k��pⱛR����SC�?n+=��>�f��-��l��М���H���X�6��RE�~���l/����g�y���+�懞���!����sœj�/���Y�]��T��(�_�'�뤴����N/r�d�'Z���ow�9����e޲Q��!5&�2l.�����E�k���e�F��`1à��0�(��B��9�	@��a.�vk#dg����ه2�j��cG��i
'�U�o���7cg�}W�����o���D^�z��&'*�a[x�>U�3���at��Ќ��J �λe&�M&l�x�zg|��7�EZvp�\��������g@�����"ۜ����$����Nlb�a�w�ӳq�À��W��p�S�w�$y��3)��f��&��~.��*��z+�?C�����P�`A��RQɥW�������`���Sr��C���=0�ݤNB���z��Z�1`g.���j�K��~��T��w�t���0dB��Y&T����׹�	�͙&���
8Ն�6�1�~��h�"�5��>C5����KS���������?A�Z���t:�u"S���w� ����[j�4����1�:����cÊ��F���X l�@��!�N�V�:�����z�ۘ�����2ղq��h�����i6���ς6R�A�3&��t�N8p0���*}�y��0)6�`�����*�x���E󉜊�ԕ�f!��I J:�֧���vl(�l"���L��/�Ĕ��*��U��P.g,�\��F�cq�{M�x^����BܒBы��IP�! N���(�p�����Y� ��q^f�k��D���DFn���5L����׹zK0ƨ�$'��;9�F]�Q����b���V8^ݭs(4����f[_�~�-xO ����fD�E�xhJ���.���N�I�v=���o��A`'ʊ��ӿn*3�[���ƚ{zBY��k�,���N��|�!��r��v:
��8�x'��R���6����8�F:�Æ>��Tw�D�Ş7��_n"�����r���M�z�� ����^W�t6�N�.�U'!��lV0���_�/󡗅vp�d50�/}�ߋ��ۓ��,_}5�/�RW7�T�j��MG�*�m�?S�>[]g�(�f� ��0җ������d�,/R�2,Л���B�=բy�#HF��3�j~��~��mj���'����"8~GB*=�g�R�s��d)��+|i���X�Af�ct��,y[.m�{�m�I;Hڠ6���n�;���゠��'�۩''UW�I2k����y�e������s��#�ɮq��Yl��]�A�]	]ZE�]��G��b}m�ږf��u�t����R1�����x������zB��z��6�vE�ܢsx�;T	/*n6�A�El͚B��
��s�b��=%�ቔ�W��5�����G,�|gӂ9 ��\����OJ�X	uy�T�˹Ǹ/�OS��^�D�kbO/�ʶ*�D;�����k>���(���Ġ����4 ���#Ӗ�%_;��(:0Zˎ���ݗŎ-�D;����`��e �U��s�%��.j&ܣ}����^ր�Y3�T�x.��݋yƯ"�(�1�f?�^��!H�-�n(����7]��� �|.�0Ҁ������g�֞{�P|����Ш���UQ�z�B��7�nt]�7��0>Y���7������E�V�5�W��A��O����m� ��65n�W����� �*f��|[o���;whQ�;PazSrN�+[u��-?�̦!2(N}�{����a���gs�lޘb�r�R��9�ߨ�F�i"�0�u���p�L]���[x���C�l���o���	�|����'�ؗ��I���[�s۔����)���W��Y�����
/*c�Ŗ;�{ 
D|��B}���?�I��Q�|�dM%ۧ���ʝ��]0/)�:]��F��G��s��p�u~;�|�0�sT5��[Ila�_.V���E�2���7c�p����%Y3����fnd�Iu�ݽ�(M��tDDuX�b���*��خ�e�l��Pej�$y����Єɩ� X)޳kRV�d��r��Jwɼ֊P/T���J����5;�}A�|ܭN��k���t�<(�U�i����.r��a�#	¿J̠�冭���<�"'NH���c���//M�6���ق1�E����i~6�CWK�_��e�0�nQ1����+�4(����ݏ����:�1��H��o8��^���-Ai���' ?�^����x��d�;�*-�c6q���^��yO�a6�,�)[�ֵu �.�D�@������`����ܳi��/!p�?o}f>�8^N¤�w.ʼh�O���f(�#��zs�
R;�)\���`���a�H���{��M���|5!�6�t�^D�����
�x���"5	�R.#?��z�zw�Zm3�X����h���� ��"d�u���ⵙ���ݢ�K�b�A�N��<?]b���)H� ^ܲ�BFeZ&t��O^hBt�@l�=S��8B���'��f�L��BU��=�	�l�i �p>6w�-�n�4B�lX
��:��i���7�?�A�Q����i�W�{V��ay!�X3���OA~��a���1^�Re�i�������Wڳʆû+�U�ޛؘu>$[y&���*d�W đ�����C���4V� f��GW�-ȫc�!$|<z���4DM����XN{��$LҖ|�^��7�?�F�0FD��}*��ru�<��ͼ�'S�i��v��ģDƍ!�����t�Ƌ���s�x$~#���0��y�~b����єq�u��o+܌/Ǽ����nz�n����,���5������:ll�߼$�фÌ�f�I��9-��ǀJ`��d�_L���k�[pg��*�7�u��.����΀9f>��gb?�GC_m%2',�$�����j�nVhs�,���y̜o� ��©��J�u�R��#QHFVp7֩������V#aI��z�����0J��=����d�	誘|{$H�IJٗ��52{+=���@�C��v��]��T5%��Y���>����!��ie^�2���ãm�
��b�Rٵ�����:L�����t����7X�X���_��4�֭;.?��X���R���e�����,�����D��L���HKsrӲ�1,�WȄM�?�k���#���s<V]"8̅v�v�~�tJTt$EY�D�k��{α��ل@�ilHQLݙiP}bh%����U�I3j�F��a���GnY9�$�۔��,��*P��Hҵ��_�6r��/���Ξ�ͦ;ƌ��\��Ǟ����ݲ)������ڔURh
��_�����W��7���/f���'�����tz�f} DG&#����N�U�b��L�ŕ3탿5q�&W��Ӟ�vh �euLT���M0�;��J2sz$����{�< �#c���"5�cR�O��l��6��+��צQx(Cș�3�������߮����5��h��b�z��k�![Z�o �O�K��,vں�U�5�����k�����������n�%t�cZ+�X��>�/���Jo�K����Ě��^��0��M�B+}^genW��E��1-��Ϟ�B�c�����:�Y��� �r�Td<�3Bh�1�%�����1'^"����S���:��t�����7���Ь�/�c��ZÙ,3Y��g'�^,b`�+��������`]a�G㖈��&~3��c���p��{�b�?�T�J��VH/�<� @����/��Re�y��\��_��L.v�|�U�CǢ�gm�{���bxȪ�e�7�?^l�Cm�+�i_�_3a	�g��I5^R��UP��]���X������sQ�?Y�/~��	�u�GQf+ �\�z1	g�+�=��z�����tz�Ц6��>���2B���w������P>�KYR�%i(��ôR��1z��%��ȑ��}ԟI�������7��"av���u��A��Ꝟ�:��o��l�:y�c<G��LcŇ�V-P�,���T�d�A׽@;)AI�����p�~.�c��������;&�c�,��%��������x+F${:Yle}�5e�P�v�6Ḍ#?e�!�c絛>�Z���	L�bXD���	1�������O	�k���Y�Ǿ�UZ�7#aĔ�T��z[{h�~���]�P<v(�$�-. 7��T,�%�qg�P�<��ȴXMFU�S��b�R�"�)�+T<��R������^�1��f]�_�~0X���K�`y�fx�ϡ����;h�5+���d�6�ɼ<"M�Wor��|<�N�㡞窮�V]�M��o7%x$i�t4���1̠�|�-㓝Ph���l��s�������)��S�euV���ٸݚ3�uܺ�>��?�����_~Aǻ�x$"H �1�]���*D<�$;��>�mT7!tW���:���9_��L�3���H8��$K�(�sw'���3���_��3��_Q_b����
Y�,��G��C_����� 
�J������6�����"�b΋@���� };[. 噗K��^�����q4�Rj�{��w�2W�!�TG�S�ȼit�dog�ӻ�Z銬#����{x�#�x�,W�`(���vU+Mh�Ais-o��7�����t�|,	pݖ3ۮ+�|�}综f@���
nRm[#j�\Vp� C�P�:Q9���^�8rv�q�;b杫g���>�:I�� X�	���/S�S�/n^�7�3K�o<�7�;@ڧs���B�\W߽�|M�p��]�;b��b7z�я:{����8(�2�f2���ſ�eH��:�!f���C�v�U}5��R����0�
l�n����kǠrk��	���޼Q�4�5��Uv;��Fu� Y���Nb6�A�;�<�;6N�E[
���|)/o�g��B	j/.�[���9��(����^��ڗ�^}|,�����y5�F9���a�2`$���^��B4xh�0t�f%���4cnY��6MK��n���-'~��ۋ�/sӾ7�q���yv���@����l�\4#tF�Fc&M��x����JU�-�d��o��y:`ϥa�3��uk�FG_��l!.#����+&���" �v��Y�^�ɤ�_:d�ı����Qu+�����t��>,D��>������솳F�~�:螘��~M%P������3bX@k�]��<�o����'x���F_����O�\��C"��h
��$x��H�� "�%tHA������$�01�%s���鞏��;�qu`3æ���pQ;M>��g��Z��~-f�|S���	~��Ȭ=�w���-�n�)@��H_�K�8�ӫYL�Y����	�O���z��L�p�Ɗ18@^�M!��r���A7����h������{ʸ-$H���C�1�LրbY���	����L����8ق"m�!;�ͭ8�@�5�Ʉ	V�?��5�����f�#?�����ו�[mw��v��j�2x�g#���u��BD�&�5����`�H��	G���s�hؗ��N�DԦ��@}��PN
T�R{m�?�EG���D�����6�q*��������?�u!;I&{H��"	�8�~X����[	�f���;|��v@^A�5Q6�yL�+��\��.�6���Y�a?��s[Fp�0�̘�׺�Ŭ5
<�jdR�y�o�I�r�w��?����KH�c�w�3��9�������<���]�"jQ±�!�v8�㕙M����d����kP�\�p �\O �G��rg=!�,֒�?������z�H���z��"�>�֎��B*��c3k'bi*�S!��'Ԇ���u����ا�t��G�Q�^�񺉴�z�('`�c|@��i�S�S�P�7^�|�%�S��+�~�\F<>���<m5��3+``}ɴ��*�o������B|��)b�:�hO��ц�Hހu���f2Q�n�(�����.�9�aD-�MI��Y�diЉ��l�Z�5^��Z��~yef�L;Hu�Z�.���%�.�%
�BS���O�>�c3�G��G�j$]���<]���a��,B�]�-^R u��=��rC�P��9ۉ��_;Gg�[#�tKnW�f��m��5�/+�A{��-6u�]�%�8u��p%m�_Kq�<Wip��^7rKj����yE�����Ss,8�Y�d5����˲��0�/�,�\![���h#e"xj����{��(�	�}!��:�q�}�p�(�z6/	O�(r�2�O�1Nh��q��pT\RO�xۋA��44���}(�I�U��s��Q�5?�����TgU"ҳ��2+�O�J�f��K�,o9��`W�+���3(�,��t�V�x9^����o>a��¨_x�3yU�Z芲�X/�db�mBH����qu���3-��.�HyO����|�G�N�NeP�O�=K:h*y>U1���EƯ L����T�Ѭ�A�H��2"�%�pm�3�^�C��n��k�s V��N�����X�ņ�Y���$X��a�p��U�V��B�	�w�tw�eȻtY��I��M\���Ӊ&���][W$'^�i�61{{\_]l|�'�8��s�)�e�6��C��~�p�߉�>;�+$�g{e��N`_)jtZ�c�a�e��P'�Z��-�O5U����*q����`*F)e3�ֽ�?t��\�W����5�����	"PD��V��M��B;٭[����}�b��Iΰ�5oBU��$F)����*Tryؙ{"+8V�^��.tf�rJ��ؿ��<|d�f�RL��SVdBJ4˙������*7!ѱ�=�JA{d�?���|���wi3Z\�(ij_�����1B�,�����Lsy~�7�l P��
 W�F����������H��T/�"!F������I������¨��]���x��wF����?�e!�M�ӡ�浽n�zD&I�	F�:w 	Ͳ��[)��q�^�\��b�B̈́��[/���6Ɍ�ʹ�	��︦{<W�EI/8�l���w���_t�2_���sX���-��a4(# p��F�����A�
~"ɯǧi�'���KPz���G��5}C��9���9�:3q�~Ɓ�8�:V/�s�f���;���h#a��q����$2������;�:�ϫ�٣e�@���z�RW��BYi�����c�b ���2�T􉭀\�g��Fv��g��غ������,f�A����5�N�������\�e ��8�W��dR�1����?�����Vk�F_ d�ݳ�lQ+����R�7����M���f鷂��� �<WK�}���n���O�Y���ϵ�����W�p��i7+Ոq)��E����K�\�@��>��`yO)T���"��x<�~cwE��є]z���9!w�[FE��@@�$��k�(����^����lN�\���V�gk
�K��1��i�%�L!����ͳ�ǖ5Q�?��� =�7*�W��M��9B£38���G�3rW�(�<_��
A�?ˮ"1��(��4推�W,���G,V���zBk���6Bq՝pS�<������z���_��X��!i;.�5��XL	����sf��-t$m���A�_b(~x8�Ѻ_n����J9�I��XGS|@��y��H.�*/���U��.?_��t�����|,��E��'pS����jø�/�v����G�m�xf�Y�i��Y�ꡛލf��⸡��Ӽ�)?8Rh�%c��!�C~�<\x��r)D���} u�"�'�gޥ��Fޚmk-Mw.ڑ<�,ejE�O������:�4�C��8V5���ؙ���+�	�87�K���(H��8���汖�e0x� )PMgi!o�,�6�2J�/>��Қe8œ��=���`�jo<[A��D��q���-igV�9ش�0'=m�0Q`.����}�E�l'����m��٩S���-s�^m[�3�'�>�+��SIy7ݺ��#�����Y:��QM��k⊈��� n�'}@㔟�%X�??0�[��u�ů���^�:�I�H��\�����o(q�t=�̒�.�O�ǁ�
�.��O�@P�,*xcq�/b@�-c�(S%��i�,Ǳ�jK2�� j�T�kF��B��?��[�-C��3�����L���dӰ*:�y���L�7�!�ov�r�96�-�������HiTB��EX�S@���Sֶ��0���>�sc��	� ��lP�u��{ ����b��R��G?>�M4�1Q�΅b�C��&�D��*
}��l%�^����Ȑio����+LQ"Jrv� ��j`�S<��̡�s�$;:
C�d�&�O%�s�Oz$��2�t����lp���E�S~�f�'�Q�٧����ax�OO7-� �M?�y�� �+<� �n5�l���P�HEqMRNnuT�l����E��l� '�[������]���tm���&�b3-o�k�@՜j��-��o�O���
;�6�ǕM�\�l�!�.�2b3�S�>TӰ����9��MP l� �x�Q��S^��4jX�y���j|���=�!�ܟr�eJpR9lK\�F�=�=^1mx�N>�N����/��yk��#��&��/K!%�K;u����=���R:*�r��0]�S�`���_KW�]\4��r���W3�x���)Ź{���N����Q4���E�,\��j=\"�kX�|�*���|ĺ��90�R�=�l\�C-]�ft�a'�N��5��-%+�G��ΫIW�>D�moS�>�Y1���i��ZٗAۗ;> Q��?�3ܰ�v������`�0~�� �Rv�NY��������9��U.�BeW(���:��2
�h�d�2h
��*8��柯��pЕ�E�
r��צ�����^f1�X��E�yoTb�<�lY��5x	tk3N����&�"�0&�x�[��I�0�	�|�#�Iy�����6ׯ?Z�#$�ќy����Sb��s��̈�Ug����{��@.��2��ҋ�	�əgKI�
Ĩݸ��b��/����m����޳�k3-y�g( �:�N?N7�:��=�f0��x\��K(�����fI��y�i�����^[��N����'}�@i[�x��w�CY͆�|�6�7���������`�nxj\�{B;)?�|���MÝU�G�b�PC ��v�8�h�`"kq�~�v_�,�sc,�Ӂ�I6�����Q|5&7AA�F�^y�2v���r�yY@{�N��4+��W2��BUU�o}�v���.9�J�-�SlF*E�}����t�"���W�m�XÓ����J�V��?��H��P���A�(��Ƿx���o/ԧS��Y<�����T��VCw�4�]�5.�e�wz���oMD٨F�gr苿YZZnA�UWc$��[W�!� r���	OfH�ނ���b�b�;p%dA۬������ӵ��W����C������%o�;"e�Pcj䀰���܁�rV�MI���&lB���<���{�yb�o1�&ɱ�r�/�`pd�Fvh��ֈ��ۚ�TJ�D3�m�W3�v�G�;�NH����Cz�]8�� ���Ɵ_G�������l����n֝^_(�l����QP�����9 <O> *?���K�Gd�45�I� ��D�g�AL����U3R��x6�
e��:x��}b4��X]6��|�$��x!�(ϑ{=���>�=0�dN��w=&���>���S���'18��C7Scv��h��mNa	��䏅y1��_�3ӹR4�n�����o�0�\9���f�G���'�?�bbOa�g�ޓ+��ϛn�.���xY!>�dZ,S�%����'���!A���j:ꢑbbҡC>м��}s���q��N��Y	�C�B/��gW�=�bG��0�[y�-�X>.��뿔���n�d�)����kvZ�R3��)_-�(�󂲨0���ײƑ��T���g]@�f�r����P�q;$�d����Py��>���6�����oUY4z.�Vh�;�tr��DkQ�C�M`1��o%��,t|������|N�h�5����p_��d�\@9�e��2�6B���(1(�8���d���-[2����V�g�^�:-f�[��������.�6d:s�Rkn��+��m��ް^:�
�'�%���-��6_9ZA��󽟆�"-^�9p����ۍ��1n.��^�9l��b�[�<Ա~4pp�ø�i�)/i=��R���9W�mؔ���M4dAk)s0�
�2�g�𐋟t"�dg	�ac0���6����՚���	eZ�)�O} .r�9A/c���r	�P���e��s��g�iH�>NNch��f��3 '9�V=�����ޅs�C�;�-y;��av�u���t�ɏ��;���^�G֩��u:�5�#hZ@F:'��Ц&C2B�X��:�7}�-]��7PP��4���~��)ml��3��Z:j��r����mI`�cGYn��>��Ҵ�F�#&@�Ho�/�$�8�վ�/�ĩ����H��Hsz\���8T�q2^�I�H��Ȧ޿�/���h�Y�] �v��x3dm1�g+j=	r����wG�J�K��0�i�׵��nB�Iw���g��a��{�踍w�]M���X����}�|$�����-v�Л��fYaBE��b'y�D�J�]���$���c��$:d�qm��ȽaM�u��Ю:N�J�\��@Í�fv��&�dQeT#2<�ygz��a����|��r�%)�S�!��=p8MC+iI��l�;��a=�pI�`�Z~Bϧ�1D��˛˙�EEh��M���L��m��u�*TwV�x�'�ӈ�?FÕ�0�ä������ZY�u�N���/���H�.ޒ�#j������IA���'ݫ�S�q˟+�2�5�j���n'����ӝV����W��hF��f3/�D��2�? G>�����G��+�n���Q���U�nf_�/�	;����_?Ϟ��EG<�0<	[&�ۀ�$��׮�
~ڤ�ղ�	l��t����b��)��J�|��yy����(�W#�:9?	`���%�f�m�%�~#�~c�x��RaP�#�kܨ����E�v��@��-o����{�P� {N~6����֧��
*N���gt���#ۢ�r�?w�5��w$U�|Oc����22rzs���(sRo�������yU{
��I��G��tu��������O��}rao.&Ui��y���j����C�暼X�ޚ��Pn�<����k)���X��b�d�=��[E[�<��Rw�݃�%�3#���4@k�R�<�U��Th�Y�؂���H���D���ߎ��u��J�G�9��n�F����\�T���&��V��+���ט���~������qb�0�ٮ����:;ͷ�YU��wXs���l p}J..b�Ag�A蠴�!��],��-�����|�x����,�jט�,c���`���9���h8�,\��T�_=x������a��VT���l�)���"�5�!�{{�ᡬ�P�>��c}�/7�%8��<y�����DP'l��DE���q�'J�#���Fy��)��T��^S�
TZ,�sc���Y
 xKP�$�xZ*��B�<>�D�~ݓ������)��e�ٞ*+��r��-�L2���aڥk��>B٭�#y��x�d�Mۄ O��;�I)s�V�N�0>���w7[{��ʸD�O�ݽJ�B��HS/2LKt�I�*Z��y�1��q�|��w֗3��U�%�	��b|,�mT�*�E�I�cU*�p]��}S�榼�j\q��k�J����^-(Zu�J���y�������G9������<�V�{y�X���	�9o�I(`^�1>���qRrvy�_�=!�`z�coq��lp��h޹8���*����5��5�}b?�[|�p��L�[wn=��qv&'vSk�I(���6�x*�L�D�"g[�=>��m�R<~;�C�/vF���eyk��v�A[.��&f&�O��Ia�f�ZBz��w��0�v��YS�w���&q�>����5y���@Y��Fy���Z׺;�̊Ӹ�zw]l'@�wOg�T�{�fq2��=%q鎿8N1�1��6���iDÛ3�MzG�Ϭ����|�"��u>�LM�c?MJ�$�\�4)�q��;���*e�ۺҪn<2 �H��J ��(��&�.S�{��8�(X��__z�+?6d�x�~?ӌoz��!e���PL�L�v���n�R\耈��������o�aq�%�=%�����=��c�4�E�rY�����������&�1�Eco⿺�1-1��#e��J_L�Z���/Q��$;�&��m�XV6Q��%/���I)'ʍ�Rs�s�+9�-�JY
h�6*��U'��{�0�y��N�h�Ѭ:H�q��g`���Ff��,��p�X=ڧQ��CWz2�w�5�sa���`����Dm�&�X,h�6�����M��ӓ u]�P��C97����u����Q֖���??���I�����4����q�z���^`�����;H��~K��Q)�Rw��!8����w �;3�*.�{3Tt�@�,�'��3�4�r�¡I���J�N7.�X�̕inp��r��yoƛu��C����}p�.?���0ɽ��9���J��x�q��<b8ed�#�n�eLka/BA��D7c�k����{�c�	@(����
��27_�\?e��>G޻A���Ux��*p>��C���$[`���N����������9��}�m�I?���)t�8��d��
��2� �`����yY?�e���w���DՕ+W����C���};���'�g��)Y��`vIP��&P;���`ȎE�3V&�9/�R�|gD\��]�\90�s2��Y��e%]�g81ڔȅpR���������C%�� ���3�o3�l�*P� ��@JQu��{���٤���8È����ǌ��(�la*~sْud���B����UO� ����v�e�(���l̆�И�K)�S��$	##~�D�o�_�7��˹����g@ĺ%ᒲ�A��i�����������hѼ���ιK��`.�k�N���: �򫖫3L{{{��}����/�񳾿��D=σҧ׺�`(��"(65�c9?qW��D��O�#�]�3A,d�HS�E�|��A�yH��˥p�V�4�u��ؿ�3f\��g�U��Z>fS����7�f̸>��(vFay8Ĳ�eIr߅�R�9�$E��uE�deA�V�#VFr	!���\�ȎȠf}�嘚H�'qZ�5��{��x�d��TA�C�`�0a�Ѵ��dK�vg��}u��0!�*H�6S
��@p�b��9J�i��͝��������C���/�~��}����߶ۻ�&��V��>�������Jw�!���r��R7O��e>�x�uK�3�vS���+c�����d�gsB������f�xS0��w����p����m[_U�łN���M)]�cq��c����=֙+��w��'d�{?��8�g�9/Z��5�;c�C`ƌ7��w8���<F��8����
�mָ�*��'�m�ycYLu�dFkBSʮjgT�ך T%Ҧ�.�ͥ N�����b2؇�80�<��1D�@Dw��������?:P��E�/5��#q��_��a�v!h�7�4�-��
Y1<)&%�{ӝ�t�O�����"�[�E۸�dIqH�����Dh�;�IC��(";J��T���b�4,��l�1SM[������'����bۜ���M$Mx��5�Ͷ�����r��ѣGT��9_�rgO��ݝ�92���i �=�)�%c�r7��_7x�;��s���f@��qe�*;��t tu�d&&���EJi�3f���c�P)ى�uU%�$����A���8S�U��2kɊxA*�u�<��b�ٓ��f�b� ��D�u��K�!�vM�p�Ѭ�?Q\-q~���%@l��0�1Y�h/&��V��B��	���!�Թ���h��>sE����$[�?<g���}ї���t�,�u����2?t�NH.U#g B���&F�n��lH��hC%gR�ڼ�˜F����!��]�F$T���>u�6�9�<*��ڶ#&>t�g̸n�֭L2�s�3av@.�8�*�ٛ�egOb�ۂbXu<v8�J��+�^g��ոu��qŭp�bY!^����#���l}VB I�W�R.GqhN��ڰX��Ͼ��kR4Z' uNs���B^@�|z�ĸ�o�|������w��+a��5|�2�K"�����sv��u�F�q>S [�ax�����7Υ(����@rO���_ڣqQ���h��\U�þQ�V�����ǑD16(���1m�c]b��Ϥ48b�n1��'��SVO��Y?n1��³>{���w��
�MC�5�o�<Z�\�)kj
���A��;�3f�������A�W�U�gХ���������2e��=�o*��<� �B�i[4n��������1�47ٸ��_`�5���iE[D^s��2,Y8��o{���}�g�rm�:=��0��	��o���:�_�	9/��HI�1�;��~�e��9WS�Ź�*=滷�����c>��K��o����#|� �T��J?ϐ��jx�c�%Nʅ�b��{��ʮv�W>8R��)�pv�����������=_|���$��Y���% ���p��?������Wl6�ݺ�O~�~���qtT��)9��o~�'������.��]r�3f���d(jYxw����R��-=����wW$ظ�v%X�z*\a=������z>�4$�5��ޗ��2�J��6E��ˁw�{6ȉ!1��͘�<qQ�֦M{�D�G�gJ������A�YA��I��,QW�6-�?�ﭠq�_�����#UXpT�
�ӖVB��P�[C��-K?���|�㏸�����.�}�$EJ���@�=����.�qM+<�	w�֧_�WG,������9���AA�ы-�/�����1�����_���=��3��7i��hUъ�h�r$޹P&��!����N��gR/�I�����p輻�o�[˵��:�2���=����r�C����������q&G$�"�R�ےڔ��'?:����/~�����7x��	���k4*��6�1���1�����wO�
��
��;p|�s���7�$K����GsO�9��T%������,e�	g���[�4~�*!R�����c:�����|�m�""������W
����x�[u���"�F�G�Չ'5����'����g?��(w\�u�1s8��T��ȝ��
%m#��]ͻdCwƷ�����N13Ek�R{��o��?���%�-�����?�l�k�񳇸��,��R4�{&z�Y{[�=��Fl���
����x���t�qX�W?y��ށ�7�&���;��/����}Vw��6���EEz���'>|��k��Oǃ{_�'?�)��������?��o����_sz�����ӟ���~ͽ�J4ˢ����ٌ�~���D����'b;�9דoh/�sY_�5ķnB�j��!fƌO�aD�R��y�^�N� ��R�g?����?�[��015 Fc���?�ѽ{Ļw99Y��ᩈ޽U��sB�(�Y�D�����3�}�G�Y��Տ����i6���?��������s�6l�K��)a�DV�g��F�I���#�#�f����鏎�O��'��n>�����|�s�6i��d�"z�vs�����}�.���?~y����o�&��g��g����gܽs�����_��_�?��?������>.�}���3f�x=Ѝ��y���>cƌ��`�BK��"-ue�V�PX�Ǜb��i�HX���3���g���wn�������em��?��j���G�p$I:�p�g��y�������?�՟���6�O���K~��;���>_?Z������Q�qv�~*1?�a]�>J'TR�}�����?�;w*�(.*w���>�������ן����H
�"T����V��1gۆj�DUYT�;�o�~����l��p�}L���
� A��ͤϤ�2cƌ���߬���b� �4������w�)_��q�.�s�����MDz�����l����c���J�/��0��s:_$9<c�
_'-�fF4�1%:c��F�h�6g�2]�:nY��?�a��*6HE�Q��Z�)AJJR�5��Dwa���ȍщFW��Pm�W���7�������������?���[���-�����<◿;�UA����&c�\b.kY��-��)e
jڶ������A������On�k8�&����	~��w��qç_���'5�dH�1��㟰:�����GOS�p��c�F���;����9Y���޿K���x�|��{8_��a��Ό3^D�`���}oC{�-Ƹ�]1�U3 }%[J��{!ߛ1�[AJs�F<�*OM�Ɣ)E�b�x��1�O��h$�^R.JɄ��=1x��T�S{�N�Xht��J>�b�E� uY$�-��	>a�C���������b|�U��&��ن�]󓯾����{~��w��ox�E��v�P�����ҫ+�P�@�&�X����#��x"퓯�g?�͟��]�O|�Ճ�O�׳Q`y�?��;���#��fM�DX.HlY.+�~�O���'�$�<z�PIŽ?>�v������bR����y���>�`r��
��J�3f̘q%<u�f�9粠�kؙ?cƌWu�+|UH��D���*�Th>�яx���G?�.����F�$K*D��V���97Sٝ����:8�8dG.I�T*pnKH����'�����#n���{_����<�Ư�����?�����w��>���?���xp��#Ղ�-޻���!;gXf
S�,j�Kĵ�y�.����G|��o�}���g��:�im���o���;�ۿ�����<|�Ɲ,I�ܸ{�w�_����������d�N����x�1w>����$x�Ѧ�a[�_|�����P��j�xp���3f<=�Z�pXn��fA:8��'ϧ��A4���x9�/�	Vl�D�b�r���Fe�����＇?;�t��ן�¶aAȎEQwޤ-V�<h~���9qQ������U�s(�su9�Z���+�L����	�G�3��?��>������du��?�n��{�P�m>|�]���1������1��?�?�����<lc.�u���\g�px����`;�����j��ж[*屮�n��~������M�.np����7E�t����h���ɇ����|����H��w?`���~���o���i�5��͆O~�)��Gw�s�i��Y��<�w����*�ꈭ�F�*~�`͸�e��NT4��*͞+�{�9��$�A��Z�R�������uH)�5_�^�n�n���~�g����?��gžn�x�U�^l��p���QKDK,���T�*>S�XWߕĹ���@��b1� ��s�`��N��aiB[�@8	<�l��t�v����{�������Õ�)�{��H�A2Gh[ay����7�h�{Ѷ���%�.�b~������ۮ�|�BUl�R�Hܞq����?��~g�k�Ta�=�������x	��8��
��GO��:�_|�����|��� n�5��ez^g�"储���yf���R�����$37�.�g���6^0m�&xod�:!��}���?%�4�X�<A�N �,�$B�Y-�񇯾���pc��ݣ%i_}��o�n q|TQo�=�b�L� .��<�������;l}"�-�f ����7�-��o�+���|X�=�I�6e��x�@H����L�8��L�B�Q-Sl����U3 �k�����l���t'�������Sf�x!Pw�@���Y���^-���\ȑ��=�7|o������f�������#��EX,+���j�{wش���\=�����/�� �ͷ� :��<�9�nI�d|����W�����{�AI�#�Q���O>����X-sɜ�B��������ٟ����x��)N*��M`��P�^/D?N�n�A{AB����̛�������9���]��ˣ[tb罈z�i|U�������#>�U8^�pv�l�B�� �C|}�Z>8[�X���_n�M��.(���L�EY�kz�f\��1�+/[��50�t�93<!BU����S�ү����`2�3�%D˳_2/	��P�|����>�~�9�*�)�$�ybL8��P|����F�Y�����O�>ca5fK~��os��;�*�'���Q�o/���MсE���]��/N�B��6��ք6:R����g��|���m4�Z�R�h�W���L[MZ�/����)��8<.�Y%[�@�~±�wt���T�I�p�������Ox�v�Kg�v���x!�B���ya�*���w������O8]oئ� ���hݒ�E�׿�=��S��O7��o�q*Z�$[��D���ļ9�bƌ���T��	���1�婦����]������?k�d�����.f�Ė����ں�Fw 	̌�`@^�}>�||�(�.��B��`7���Vխ�������΃�������gDdFd�_$2��mQ3���?�,�LrB���9��_�T\0�J8J�b2�(�)5ei��0R2��9_.Ȧ��e,��*��g'�bʋ����X�%j(��G@R �y꓏�b��T��W����1�V��0�R.WH��,-J���V�$y>Ő���e5���4�\5��.�.7\��=�I	����J5�zڛ�Ւqk�k6�a�Ţ�W��?��e�)��2r
�,�
%$��(
��9��TEu�����S�Ҩ�03g
��dҿ�Ea��_}��?�!�K�Y!Ӈ�)��Wu���nz�Ѩ6bĈ-��U*�9�R�e�����+rYcJ�5H�����������*��hVՒ���֢�d�22=A�{Q�,,.ΰ��Y�e�i��u�+�	
'(�d1-�f��xQ����B�����;�X)�X��-��j7oG���E�S����N���}ɺ~�R�\��b�$;`��)��ggϱ�
!UYQ˪\rp�SUp���}dv��܅��pv��
�<�D�!�X�5X�dzⳖ��m�1}�r4�׃V܇h���H�-�OM�CH��VN���X���!�:��H�Qh��h*pT�3�9ǔ_P,ϸ�X�,V,�t�t:erpH6=��	:?$�P0��)
�bU!�)��)��P�@TH	ز&o�x�Xї�#F�v!��D(�Z�*����Hqid�j\�9\ ����7��BrU��CGV���d�e���o���%g/�����Tq0�0ɦ�=?�(*.
CY9�������{�}���brx�ͦ\�V:Jgj�Ġ�u�'��ڷ� w������@S����9��ʞS>��/?��/~�sΟ=F+MUU^��V0`V���1ӣ��}��~�;�}�ûr?��O+WQ�JPBH�\S�$>vǈTIJ�ٛ|�(ŭ��V:,��TM�7|̓w�a� ώf��Sqgv@f`yq�ٳǘ�)��G<{�����1g�-Ω�K0����錻�~��w?$�����L�0=���4.�,�rE�J��dZB�0��̶a�F�я+��W�$�5�
ky	ʈ���ޟM	&:�*_@yƁ���9ՋG�ϿD,���g����g��O8�%��sXaYUe)��4P���E�ٻ��<@Ύ������r����st�3�,�r���%N�+�"�$!C��- ��C�[��J�rK����>���������o��ٗ��cQ�M�ǅ�j��c:J�p��,����'�~qBvp��~��9|�w��&�ɻ�;|�����x��Y��|,#d��+R�l����M+��	h��k~�����WW˂\:2��)�^<���O��?����ї����%���ea.B�6@�o5vi�����=;����6}�<x� ���LU�i�#%Rg`����Q|��ֈ#�c�J�`���x{m�#^�"���i�l���g�q�g�J�l���/X~�{�ӯ9���}��xJN��4�;�P"cU-AI2�ky\�.p6���H���ճO��߰4�Cv��o�������������R�	��X�.��j��3+o�	&��dQE�b�r�-��3N�)_�����٣O��rw���3�tXZ�T��t���%P�����#~��38�Kv�~�w�����y��s�T����*����B�s[��%����N�r�.?>��C�Ys-�@C�J2s��:�?��|����׿��=F(��5�љ������IﱰeM��J��%%��y��ǼX<��'���7���7��:z���z�S�Ee��>�Q�EH��<�%�ˈ7�.Ě�}i���W���7���C����<�I�>cH���!�{�/[s}���9bĮ�g�ܓr�DLщ�143�|X7�Oj�i�:{���oy��_����q�5�\0�9��C:�k8���T�)�d�Cʲ�.&}�9;�`�\��lA�NY,�x��/�����Ï~̇?��y��5������`]+�N���ZN��t�
wˍ!��i����(��IRQY���e�J��1���1_�O�#��cԋg�s�N�H��i��*��b*4�
��0���R�-��r�*(J���1��c�g��>��W|����G�x|�$�N(�7�;[�l��S�'q�h9�zk}�d�Rxn��q��/����`>;`Y,�+�\:����G����Q}�+0��Ls89�3��Q���- �q��!��ˬ��낺�(�ݩ��V�=�_�}���o��������!w��yv�vS��Q)M)��Q:���sF�=���a#F�
���:F'.K��Ҧ�B!�9>�:����]����H���9��h�
�*��u�Ɇ�.k���)#u���8���L	�\��g\|�3���/��7��^�`.�-����uR��T>���>%�B ��?�V�͘d����<{A�*X+�����9�x�����������>��
���,/��3�7��g���rE&JՊ������%���d�G��ϙ�S�p>��@�)��o%E�N�,dJ!g��,�T����ł�r����O~�����+���s��!/V�lJ�Z�Ł'��H��A 
�܃�C�PdR2gI��w|����?b���s��M�LU��|�l��2M�$R��̦S&��X*SQ95=�9� e�ʔ�y0�t��E����������������R>Q��q:�.B"�/`(�:{݈7/��ĊQ(�,�*�u@
����mb@�}S�z�*R�pq�`e孷B�8��@ܳ�x��_��Q/>��T0�-Jd�(MAQ.�2m�U
�L�R�_�Z�1^��X,ȴ�:���M�YV�a�\�b������:e��k����)r�>Fk�4�|U �h���1o�#ݶ~�`.R_�ο�z�)����^|�K��)+��l���n<Q1T��Z��X\��y箙dY���I�$WL3��rA��Y>��_�����O�������bNiP j�X6���G�x�:��gƲ	8IQU���s�g��o���������kt.���u�a6!G2��L&N
LePRRV^��3OcsT>U��/� �͹X,�f9�Eg_�����g|�O����6���a�c%h�u����m<9bLu=bĈR@ސ��zo&q�n�Ǩ���e'l��G���^�����ӟ��W����+N�W�KK�\�O4R�4��N�����$��b�����}6��Z��JQ��%Bfh�'FX����|��+��������7x�Zal	�	�1oC��Hl֚
�*��3�x��������/��������*�J��uLG�ЙFIEY���,��}��j�1�u���t�vyN��|�W�3Z
��w��h}�p�V���,�o�K$�I�"��VdvA��c~���{���Er��%�,c:��*#���T(]S�E]D�,�K
�)���Xk}6����0UEY�L&�H-�	�����������������RAa}����b]��S3ߌ>1b��c���'k��1F)��|�~�:UU5�Ƙ�G*�����M�&�#�1^@�u�N�I��2��B]S�k(6\G�+������[�L�	�KpKT����~�?��!�>�n�d&,��~B�u�9�$? [���8Ge*�3X["�b6�Ba�R�\,ɴf�Za��:담	������,�Op���?p8;��LD��&,+PR��tr��r�n^�P.���;-,��)8:�����3�=��/��s���xx�;��56��^M��,��m��Z��%eY�eYK�΢3MUV�y�1�\+��2�4�f-(�S��O�����T|���qr�#�]X$J
_�0��m1��S�[����I�9;�݃��������s���D,s�f�d��c�����Dk���,h�)�r� �aJ����+�������H� L�)��9�\Y,8��o��{�w�P)ũ-( t�y�+���b���q�k]\��l�NëF�S�hD��u��F:�կ�9#F�k,EQ2ך;*��������a���;c�C5A�)�j�H�+�MfŒ�T��e��i���<ǖ�i�,k� ��_�\�Ȅd6��WJ���g��_���Lr�?#;z�eBU�P�Z���N�d�:c�
�>�-����b��7�'�@TL�cB!������:�l:�(
��UY5��TPZᜡ�VT�@+���<���wX�fdg��9��ϱ�~�W��7�G��?�?0��Ү˹���!k��^�L�s���t���?�w����7�;����+A�%2��@;I�B�6�I�=���/�K%}R)��r_k�:lYQ��)�+��Z��RY.�Mfay��s>���e2�3��OXI�U�P�:��cT>F��c�%!��!5���T�qJW�r�),�o#F�8I6��ʊYa8��c>������+�����@8��kJ�Ӧ��QYS��0��J��Y>��(�/I����e��DX@-��3�	�T8%�Y��N�e�2��k�ǖ��o�?9<�drtƪ��r�V(AAp	�ł��?��	����Z2��<sHc�b�Eb ) JJ��(kq�a*��)%��sWa�@�j�Vi/�j%�&��(*�̬�.�����K���;�}��7���ަ|����T__��,X���q�.��Tu6^�iDU�%f�O�����?����p2%�5�|���(����I�]�p�#��;��S˳�>N1�(��
�T
)Af�`i�؊Y~HY��Ͽ�ӟ��{��P��X:O-oH��#F\=����\]+P�l��|����7~��\6N�Sz���X\�lɁ9㳿�s^|�k�T��L�1g|�:�VhU�:�3�gϞa*C���yNU��y�����9UYb�EI�T��d��k-e�BX���J�g9�ٌ�4'W.ÓO����=�\���w�`��7	!��ׅg�vŬ:���?��o��<��Q��,GZ������kl�|8��Y�� �Uټ��t�I�^�YY+�Z_��8�bu�҂Y�q4ϙϧU����|���@�>b�A9�3���a-i2������6�����,.ΡX�p*8��g|�����+rePY�Χ�,#�s$¿����)X�O�W�'�,;稌�,+V��咋ł*��9V����4�v��3T���ͣO~��,�\��DR�U�)o�x]��ߝ���|���xX��э�8����9��:n44�����TX�RW�7����j�T	�,vbR��n��'��Ze��Y�T>i��n�&�֛��p��hB8�@Y�szĈ��ˤ��4!,�V�Z�(��L���-y��?��o��#]0�q��@I��Pg-+��,���>�0NR�
_�BH��8_,�:Cj�ԚE��ZKQ����s�b+��x�s8��:G�eb%��]<���_�|�;N�2�������P��kO��5����c!O*�5��[�ʕW��L�BڂC���gT���ܟ.8�*�8#A(*�pN���Z�g�9���''�,�8��t����d����Aj�u=�ٱ�1�{%�/�
��0�RY8:<ƼXQ�ͳ��%�?�!w�{�|�O��E���V1L�����SC_SƦ�;;���t��y�=ӊ�� {�{����)��|��pY����t����+g�H�V�����H	�Rj���P���TLg�V�f�Z���D�|�mk�l�T�`%Z�1%JHІC-���?E��q�����/��.~��ze;FN���c�nz�U=�l0���,|��{����ZAY���X�:�����w�'��Y��k����n4YW�~��+Y6eG���ی0���):ʏ�W+,���ČaE-�9o���U��F�mH��{���1օ�,SiY<���_���<�h�g>A�p�u�u�UH:�����c�O�v�6)pRQT%*W��`�X-Y��O��m!R 3��2��L�]P<��O�oq����
[-{<��	�����,���_Q>�-��c��I^��W0/��*�(*�{CS'�[
�Tk:�9����5?�h$�@)�V�y�3�Mɲ	-QfE�����_R�~A�8Ô+$�������W���kE*gɬEK8����/>��?�j�d�1;8���-�g�(Jt��Z�b�Z5�:���s�TJ���a��Pu����3��K*2�e�x��W�gu�%J�����kV>F��^y4NW�����\Pbhd6�7��ֆ� ���~��+��=!o�� ��38$��2�vk-�Z�o�Gj��3����vϬ9C�����n����]6~F\6�n�q�n���{�G���>^�L�����B�D9=��/?�5�l��`�%VJ�!GF�>�.賳3��y�9D!��Y� �L-��EQ��%=O=�7Y�QRI�Өܠ�,*���<�ſ���~���C�9E]�M����KgQdu��_��g_�a^0�+�L���	�ش�r��8j_J�P���Zs�9�����­s��t�V'-y6�La�ȹX�(O���'����>�x����}�T�bYg��5�2޾����SԊ��"�D9��l���O��/��}��4�,�"������;��0f:��
����UC�*˲a3�EI���*��Te� r�"1|R�֚�:�8���'ܹx������N���׌��G���bh筗��v� |���ǂ��[����H@��Z6��a��0�|��V��W��mW6�X�_���|��L�D�c�u^�
՝�;�:�����c|���d�t:%���K�,��J/�@k��2�-�\<����J�|u�7��dQ��x񈧟���ǟ+�usk}��<��t�ޢ����|��u��DV{@�c��X y���/.YE�g)�}'�	Y��2nO>���'H��٥�~D1��W��.l��.���|j��j�ٓ/9{��1X�t:�����K����L���t�R�,��Z7��,��S���:�����ł�b١Y[����g��	ʔ�hj1�'<�ⷸ����y�X�pĈ[�����w����:bJ���jN_-z
����	��<�YZ��p}��P$��v�}�������Ჱ3n����56�}�c���&�D��9��9O��"Y<���/Gnϙ�
go�����N��_\���xk,��(�m�PJ#��,��(�%ZK�R8������Uբ����V`� �3�jB!P�,�ŗ�!��:�Ybo8�y��!�>
J�v�LV,�c.cW/�X�-q���5+�4EQ����l��GY����:]oP�U]T��A������fY�����/��o�RZ3��X,.X�S�}��=�����D�r�,
mZ���^כN�sI�b��/���WHiqՒ���Y��lE�ZB�\0�L���?��9N3��0eI��_�
�U���!�|�љ�Qm��,p֑�x�x�T��rI)1�i�[�Y�R�|��ճ�X<�����I��q_�b�/F�>�������&�>���z��놵�@!ĕ�?A&�Rru�^5�(X�b��.n�2�����o�b�c�Yx��!j0v���֟��L�a*�L0ӚҬ�Z#�W2�М_\PY��tJaU�.TH�d���_�����@�*ʂ�2�gM��]��k��:V�����CW�Y����9e�|�K5@X���,�a������L�F����,�F0�:Øʿg�T,X��}л���ቡ�$�s���Ȳ���	���V+*�PJ��Bʜժ$��I�\������,N�1{WP"�ik�tk������H,Uq��.�.f���b��%a��	�@U(���`�
�eXc||�֝�[W��Z7��1��F�R�����0	1�^��^� �>�m�7/1bīǍ�r[�� )��SEF���&�ߦ�+�w�,��@���L���֧��7�T��`X��S*����:�R���dBU��i�+/,yz�����R��Y��%�Ě:�V��LrM�)
�@T`/`�ų'<�1�t��L��
%�,y��ל?Ɖ��IX.�&�]�V+��V��V�U�n7��:�Ö!ͮ��B�~�.�V9Rj��}ha"�G��'�LIV�nye�V�W>�4�®3��M��*��&%d�Ê&`Y.�(�3�.p�hZ�Q��6*ӊ�s�Q�vLT�6�����X	

@UVm��t�R�xq������+-Vjp�n/qĈovQ@6$�~�%$X�,vwe���&[��xy��Ux.s�����~�6lz?W־:z��m��咢X��c�S	�m�L&�,����|�����Yʪ���jn�j�B�Ɓ�����Y�T> V�P,������ K.5ZH�t �����9R^w&��s�"�gO�.���)��Fʲ���Ɠ�eY�r.�s-��j�BiE�ed*kҽ[R�%J)��\U>8Z+�G�z���$c�X1Ղy��R`����o��jh}
	ҿ�%���[,�8WB��M��l2�H���I����@S�3(������B�A�����ui�5+.8�N���dZ*�W+ʳ�hk=uL�k����(v#�fX����<%���꽳%��o+���vV0������GD�
����>3Vw`:��V�Z0��Y��{�|��;�p&_��f�`a����n�����3�N��ͩܥ?�&t8�o��=��>�5��|������&�v(YQ;��`JZ�+XU�<{��aU-=�*R��r�k��L{+���Y[�hZO�V��1���Ȥ�(RIr���d|j`aN��
�W6�/\�Or2�P֧�u8����g�_<B�ᶦ⽹���ca/�Ɛο[W8*��9�\p�%9�=�(��2&�	��k��p�e�&�*O�5Vsk+��)eYԵ%,��:!!�T��MJy�h�_�Ʉ�,��
�g�Ϲ8}���*�PI�}�u��X1��k����k�a_������3V���,�g�x�� Ag
'B)�RX��J���	-
���l�ύ5,���)uZ!�$��5]�U�LĘN�d���Jf�	��|��	0=|�-��pv�������/w�֩�^� %������|���y�ͪ���_^�_�X��K�%���p �C���+����M�Ɂ���bp���|�*2F����A����;ne+���6IR�N���*�ն�b+�Ul8>��$�����{�����YݲNƤ���ug�`�\zOG��qm�,�JH0.�P��.�K�O!�R\!��tLg�b@���1h����\	��7$Bʺ��=��\U:�	4�d$��������Eᕈ�.d>�k�=Q����ZWX�R�E_=uSbm��������vj�P��F�i~wZ��3���J�l�p����Y�g���s�z�΂e�AI��h���y�.���dJd�5)8??G��m�JGQM%���WQ�,UQ�v�ʇ�_�6�fĈ}�.z
���dm��_	qsc@n�T8'�&�v���P�؛���R=����:�j����:?�S,���T���V+��sɧ�ioV�4:X�CA�ed��c�h�׃�|>��!AM��Ae3�,��W�D�JG�k����0Ʈ�9GYH���K�Ѻ�r�\g��{-"J\��bQ r@���cZkt��~����TR+d�#�"���`}��U�o�Ĉ����Y�~��s��IQ�1�k2����x/��	
B�iy-F�y��U���PN!�h�Ǩ��V��ux�X@����R� ��d��&��|ݏP���W#F�������/���)mNlH&�p�.�>�`b�-봪
!2��9>>����l�u�����r�P[k���5��+9��ֶ���`���,X�c��g5-�IP�	zrz��a�}հ��*��JJYQ�2�M|,���e�d�*�`�@u�ԅ؀8FAJ١TUUEUU`*O�2�0�N�j�}�W�TS��X0V�2P�v��&�mP
%�v�f�K�H�>�M].�>Gg>e�Xϙ��H�O�2�N�Wʭ�W�4�,�F��N�����s^a��:VHBa��	B�,e#F�ч�
H����!����q1�~�4��ebU:�s~�"7���lc�iG�@ �����N�Mb­9�Wl&��Q�ҫ�yH�f/��*��?�H�U���~��(�%���� ���L󪱘��vQ�%Z��#1�L�Ck�N��r��Ҷ�#x8����-�����ҳ������YU{4�3��be�>�!��d�K,��*�e�:Ș�'X[54�u�]���W`kj��X���X,e2�ɡ½�z��9Zk�����T�EQ`���"��,_Ӥ4��!��;�L�5���M�v���؏�<ˡN��uWBb�P �����&�r�H!)K�@,����/��,��� ��c�����?�N���E��Z�t�ڴ-%&�ѓ)��#�tF!B:�#F\%bod�S���6�}�z@Fl��y�벬�	M���z1�֡��)�F�5U$�4>C�?�*��,��F���H\�<5"�X$��q�� (i��UX)�1��|�P`$�BO0V�nx����	@
��(�!�C
\��<��m��YGe����	4J_��(��+&ka��u`�W~|[�1�eI�,��<|�}~����"d��%|�&1@����c��2]���"��y���^"�|2o��-��F�0��L&�:槪�V���|�zE��G�)t��``SR�,-�s�Y:*9VB1b��1 W�P����A�����#d��
��%}��T��}X����ڒ{+��]�jL����E�A��qA�Ԭ�d�����zLe�K�r&�����y���Zd��l�\i���`Y�V�lS���>h�6i#��r�!��*Kl�s�R�3�Z᪪j����*�=$��n��Vf�&�s..�)�c��#>����Ύx^��O�r�b�(�:J�`C��+��88<`:��T��c���8�$X>�yT+'��\V���#R�ރX���ٲ��*��c���2�q~~�̟��g��a��+�J!���r��:Gꬎ��7{~�1��K%��y�+D��ĩRo�KlĈm��C�%M�&=��)NHa|�QW�4� �oG���U��1�y^�t�M��Oݫ�O(Z�Z��G��W\Ϙ�f���PY�q��L��gvt�Oak�-<�8�M�u�-�u8�39���V�s.V�Y>A״<GY'�p(Do
8��ZO�Q
�y��&
�5k�ψ��@8�:���Rb��T���)��=NK���E��'�����;�����~&����]Ϗ|����Ae-���sH�#C�P͸_���R2�M�8�`�Z1�͚;�����?�5�'1̿�d����7��"ψRh����"�fs&'w�DrC�d�[���4�}G�\Hg�^���Opބ�`�[��5C����(���ө������|5�CJ�P|K���\x�J���9�۾�:*9�/��5��Tg�`nwW�Q�g���S��S�Ɏ�������2S3)��
aeQ��X0��Ȳ����F)˲�� O�
�eY6�������ӌF�-!T�I�#gg|���d:�ً��V(�f0����K6;deJ,S�K7{=�k��e<k��(=�<���<���X=��3$�!S��X��]s�����3�u���y���ы��K�:~C+M�g���QV%����Я���u{�U�3���Bprt���1��ӋĄ2����!���jf�����qI��V6y�i�G�H���0���O��Np�)�qR(&�)���W�k�q�X�����
����|�d��:�Q�)^B8�^�y��W m��cv����	�w���9d'�G�X�#4"Z7.���Y1b������ڙ����W��|��1EH�mт����M�Q�@+����pW�Q�84bčF����8��LN���]�r�ii�\d	���!<��(ލ�ǀ,�R�w�\R�Պ�����8??o�k[Ss3��rIUV���;ܽ{�/^���c���I��}���1���ʩ��KY��1b�>yqx19`UV>[Qב�9z���K��PJbk�X������W��*+��`�\P�U��u2�41>e�jhX�2��5��X�3���	����OA� �����ӻ�ϙ���
�WU��e!�h��
��o2�����p���:*LeX.V��9�T���5�9ZVe<�eU6�.P���2�-S�8!�-2Lᕛ��ﱬ�LNb�C��k���N�<�m���`v���e��"5�a�y�Ҩ"��[ �A��6�ͅ ��;���y�*(���4"�4Bg���b:�6���	���4 V�d�
	˪D+�Tھs�<`�X��O���VT	�p�o!N�xi)�z���F���S�&'����X���/���%Z�kM��k9h���|�>��,�&N'N��¬+�+�ȳ�4�bAe��w�Am�.l�҂���0��|��<y���h��;�}�;�d��bEQ��"�vT�HY!1�Tٔ;�~��w?9%��W�W��be�L1JQXG6�5��d2�����rY{�}J�P��,�FAt�aݚ���w��1x����ǖ�U���	*�83�*?dz� �c�Q�P0X�1bD���^�=g-1�ͅ�bY2=�G~�_���:�rX!��Q�V�V7��F���(��� M0l��(˒�lֲ��j꡸��tCE;�s���1���/��w��JA� 5!{��~���!�'� ��M��H�����˓߼���S�Vw�(m�j�`U>���
���)�I�R����F	���3�T�\5JGY�M�,�:�l���Z�D��`����q��]�?;�/��lapb��8|�m���Y�5Q�"}#d�Nس6$��E����?���.α�P�b�d6Yr��}����SP+��p��,X8oa�R`�u!�A/��!w|h1�-�s�û'��*��y�*;@��Wi���%�w��#F��T@���Z���Ƿ>߶�����q��;΢��l.�e:�Sah�X���R_'$Tٗ�QF.�<C1=����^׻,B�(�Y����$JNГ����?����xq����V�U�c�S��\\\�JϬ3[�f�������k{�eh����pڛ@��5����c����o��~�3V�����������qV(,�U>������S4��}�����/}��޹�q|����t9�D�����Ȳ���r�?WE�����Z��N怯i!$(%������cJN��w���淿���8���{<��?#�m�\:��C���s�;$6� �������?���gPU g��h!�w������r峖��y�2�e�5k�p�)��B*O��כ��;�|0������\�������4�G�;1��?�\���_��5�.6Y��ڽ#.k��t�ԛ&�a��v��5CH�d�3���&�
X�=�����g��qƜ��Q:Y+(��W7������ʈR�E���� <���)}���`~�'�|�/~��:���ýos����o��ӻX48�3���<O�p�(�>��7�z�^��/�����w|!;�3�M'B:��%�� uL���eUR�EC��1�Y���	Le�⑋ł�j�t2�޽d2痿�-���3
4�����~����-V�Vz�g�Z����ʇHo�/�#g�����8~�X�[qq������X�xp�!'G�^����:CU]�w2���y��88�����-�j*�s�:f��k�f��|���O��s&����f���#���"44;�l�3bĈ�1b�k�C��xa$��wy�G���~ȣR�li���M}F��r�d�
B*Ъ��WUU!dJ���\������RI�����O������O�z�,���{��������{�È)�I��d��|X��mM�q�g�*�f��#���q��wx����WO9_�^'	¬�擙N�kt��ޘ��Ϧd]�s��&F.�R>�{+�"�?�%����X�Cf�~�?���w�}V�#gu6�$���}��8$����e��?��������ީ�-���O����_�*���qS��Y��[�=(-PZ ��J�08�K��,�Sd��0�����>����O��ũcz���w>DL�DR�:�E5#1b�F��oїG�̎�}�9��x���c��$�R,.��������W�������s�Xr��,������g�N�b@DHq-i��(�9�EQ4���.���*�����|���<z��eQQ�9?���a��O���?C��&���,�Ղэ���D��Ci�)&������;~�WO���W/����0���8�Y�*�8���1��1u�]�4*��G�3����,J*���X�V,Wg�U]1�2�L��X��g���W�0�c�f��7���?�;��|�ev�
2^����c�e[ZS�|QO�ͱ�$Y�pB�4���y���ӧ�슲x�D���S��Aj�{���9eY�X,��9��*�=�Y���LY:�(�0t��EQԵv,�C2�s��}D>�_<�I�!�}s�!��=V�!�TP���t�U�oY���	ݵ�{���S�
��Ә�a�
���I)�H#q�c<������*�W�5e�uΧ)�l"u0��'�y^l}_30@/�w��ǥ��%�2�ۭ`�@�\rsu!�x�$�~�~Wq�;!$�$W3�E�`·��;����~�����'|��%AgSd�|���d�*�V>-oY d�[�HRBeL�aN ���*OG UF>����3O�Z��\�,,���Çp����H�ޏѓ�,�d�#�}�lL��vg�k�M/��|�1pf
|5��=�����G_r������2��x~�0E�d�\�uV+�Χ��W��J)Ȧ�K*Sb�8�0��p��/����3N��������O�O~��G1.C���V<T{z�]*����K��O�H,y�3�u����������:�g����ri���z���`F�O8Њ'��Z�t�ZK�N/�r�P>|�&uu��g٪J �ΰơtR�e��lZS�,�|����7����=��31��)'�(�	i�K
�O߻����;�FԲ��z����1�?�ݐ}���=��ܳ����NP��|!X���^�+��[���p�6��KBy)H��	Ύ��2��^Ra�9�Hk� ��"�Ç?�O���OW������@q|2��h��
�Vh)��[Le8+�l�|�:ݑRsLY`��9Ae+T6�0O�^P.K���1�
#$NN���'�m���?e���QGqv�+<	��u͞m���E���pR�b�F�#�~�ϸ8=��7+>yt��r�Zppt�aq��);��j���߸�yYVa �s��D�kT�svv��ǧ<~��f�=�?���>��[p��� $�e�/��n����С�E�$C� �%��Qw��X�q��m��䌢�(d�]�S}�:�ރ�S>|�j���j�c�CjA��vӵ�2�}͝��0�"� V*J����==�E�s��������o����#����z�Y/�6����s5b_\���*оvv�+u!Ԟ+�u%t�&�j��
��1pS��2bĈ��%��_'���@!�lY1�4�J�g x���i�o�M���G<9��c��D2�4�|�sk�^ղ���E��c,ei���*+��)E��,8?;�C�2 rr����6���'{����4�Yd������K
r��X!0V@>������;Jr�ۿ槟>���y7��\�S+�u(�Y�%
��J��YB��V�#\N�k=e�I����?;���	�C����?��9��c�''�� �A
y땎��C�А����r��엿��e�O�=aU�3?�q||�Њ��AQUT��e`p>��$���VT��'�G�XË�|������{�����~�*;������ʉ����[���],8MM>�W���ZM�,q"��0���s�腳!^.�ZpYo7�M�M���t�J�B��J�X�e�ϙ���,�dr����5O>�_?��ǲ�d�9���B�L����g���UQ`Xk���buAi�LXN�Р'pp�����G?��m����=x����T���9oq6���.XBf�'�����������O~ɧ����`6�L�X���H���<˱u�+K�l8��S��E�Le(
��X�_�(�)��;}�#�����7��r���A�Jb!�C�h�t�v�*����˃��)RY>��!�O�N�pZX8_����ً��?b>?�`~�S�Z��>]U��JQӆ%��3 D>AbX����RdG��G<��0w?���PV~�
?��px�K��}3b\f��tCӒt�Y�J���t�2�C�����7��U�R�]�a�c���ҝ��#�!\k@�k���`�!r��z-��ҥ�	�A��#�d���V�1�c�\C����.<M�H�u�|���}�w�����7�w�᫏����x������,C�s�S/�΢�������a,Ū�m�x*��Ýw�������������}�>��C�ʑ>�s �yn򛷤m��
�J�3H������.jz�;KS}�[<�����kVOǢ*P�d�%�UdJ�e�B.���YM��zó,�,�s�
p�	�y}�}���[?!����RP���G�V0zUo�p��r��UL����T~������?��� F�W���|�����l泑�����g2�J�8N��Ҳ2��X�b�]%�*�;����0�����.��RQ�	Rht���:��s��+�r+��m�l�}���۞pv��𲠭�z;�}�:�x������MU".�]= o�r�?�Qk����.b�{8�M���o�m��1w=��	05m�pB�Xa��Lߟ��;s|�=^|�����)��X�Z.U�*`*(%1�]
�q�$� a����ٽoq��q�;�E�}w��J!�!r$>ͩ�׏�a-��깺���A0��<�&������P|��,?�O��+ο��UQ�u�Haj��z��ײ౪��U�)r��9x�-�~�c����΍���;�8#�=��۲!Y!1�:��������ٽ{���C�G�r��g��k�Xa(�(d��9X�+�K�T����|�+(*Ù����������G��?���#ﳲ9@#u�qpyZU}�p&ހ��C���v�-D��׷��C?��^�Ѽ~E�$3�i����>ܐE��H��+^��@Ӫ�F�A�3�@"�΢rE����{L?����3���|��oy��oϾ��=�����!�q�J�)��`$ 3O�:<����>�������"ODv��Z�h�{l-脢oR��2{�7���aa$u�[(��C�#��9'���������Ox�����_P��8����J�����qwȎ��H~�=�|�����Oާ��H
W�S�Y�\Uo/�@|��0^�=�~>�5�s�${O����գ/1�O9���<��W�'�a��%`�Y%�Z�B�T�f��'d����.w>�.��w9y�C8|��:��C���e3�ʢ�BI�uET�0�c����VOոս%x����Ԑ��3��~��W�p������\!�3�&o͟��ۖ59Xɜ�|��cp��5ܥ�^���Ijţg%m��ֿ��,m��WL��X!�ƨCF�2����?��ߧ��c�>��㧸�D����l���$.�cTƽ�?�����{����P�FL�j"�8��L���,m�c���.l�O	�~m����(��rSU��9��=�{w�����q��S^<���_��V�����t�d2A�3�}�m��m����wyQilvȩ�C���tr�VS��&�Y��$"U��i=�	j.�STH�ґ�'ȣ���=�]p��r�޷x��ǜ?���,���0U�+���Ԡ$d9�������p��oa�1�#
�qnV��k�T+r5A!0�� �Q0�A k�{����U�O�?߭�w�`�9��
����x�d!�pkY΢��Ԍ���R�}������W&#=��)2C1 o��{+֝���  �Ӄ:W��|�Nx�	F�(�?d���i]s�T����:�)���##p�!�z���
���loV$�yƭ]�V�u�����3���١��+��iPo+@Wg�Z�K�N�t`k[�c\@)H�VbE�Ugr��#O���MNL�{�"*���mA��{*k�bFEF6=1�P9�+Vzo�1gKP
'��Ip
e�mn6�d>�XCq�T�ݤ��O\vv�4߭�/�������ٚK	p�:e�!�N"�]s�HN:��r!��9��%��}�����w�8)ϡ,��a��\/�:�P
!s�S*�aDƹ�Lf�������k��p�&��x�B��z��>���O�Jb�I+QG$���7%����Y����%�8��b��N��9����\a��\Q�~Eu~���)��eU2��8<<D!�����
#$���ΰv��B(��(�������U3�6k�Z߂r�Ҹ�4�C׿��CF29�0�rϿmt�����L3������Ab�xPM�+�E5k�Ê����	,�
�zm�Tֻۭ��al�ϩ�E��Z��"�����XC1�q�]q�Y�F�% B<Q��QV�:3�uc8KV2y�ŢY6/0W�-��b����`���b�b�u����)���|���>&�������[`��I_Ȯr��,�!�
�O�*�c]-[��~�&�8E�!s���A:Dߡp>ˏ�P�$l�a]`�j�n;�����ۯ'��NLX]b�Ʊ��^�=������$_xe@H��3__EOTQ"�֬�U��,�ͫ�@�5B|�K$Y�O
�$U��H|J�Z�n=�t�s��g�a#�{I��&!Xd���
�$�y��P9B�Q�w0��yYa�'���V�%�1H)�Z#�Ĩ�1��+׊n�o9�
-u�HH���7��m���k�m��Y�^��W^�N�%��75�k��F*y�[��"���P+�W+���ai�#<��rH�r�
���uk�؝�W<8�t�t y ږC:k�[2����a��5�a�	ʶ��d�H��]5����CUKw� ׂe��\#�@8���#!��w�t!*Xϣ��	��C��V�/j�U��ye�~�t,��|H���F�Aw���_!dm��ݪC����d�����ÄnR���Z����} !���V����	E��@���`J�8�ٰ�>�)@�5D��V@�Ǔ=Vq��(f�r6aS[��E��>N�e>�8Y�� & �["�EL��#�{܍sX$JJ���V\lb8SR�TR�|/�m�c7����{�:����W�/�����_��_c�Y�L�"�s{��xq�T��F�
�K �!z� �e��t]ygh2vc=V�Y�*ۤO7�m���1<�'�^e"�R��rD�������Ȳ�pi��9����۵�Ռ/�T�B6�����	I�i�
'�X�Q 묆��E�i� �߻穔�70���>
�����������F�F��F�*����R���3�~�r�YH�jV"�$S�V� '}65�pN��؆��+wׄP���q��W�f=w����`���6�1i��:*���aFԙ�9a45Ǹ>��>c����-�P]��W�"K�V~p���y�bq�x=��D��O�Kd�v=�����V�M�]`��Qjm!
2�u]�O*�t�d�S&ߧ�Hd5�P��]�1�'��SeBmܲ�D[vѬ7-rVtۘ^�Yצ 9������v��K(2�i�������@�������Śf�
��IR����B�&;v�o���E)@H?�,xK}]T/�SF�d�>��=c؅s�x����L?[�l8{����]A	�5�'l: L�\��ŏ� ɮg����t��Y����T�k��X﹪�=b�H��f�i�Zi��0��ݿ]��ž�_���_����
�Vmc���VZ\OK���u�pμN6W+j��!�|J���1�z��Ơ�q���:��`����À������+;�2���r�|b�:��� ��8��R��<��puM[���GԞ���$�#}��yl�Nۘ-��B���C�\VG= {�9W[hC6W/���VeURV��_9ZU:���z
�VŻH8����¨��1>��m)���Z�+�p�ɖ�pY[��}|WQ�w�:бɤ��f�k�X+.�����%)�;]cl���}�Rێε���dd�3��snMaH[�dݑ�����6�P Wa�R>�'��z�d[8t�F`j%+
�7済&�������M����d�Ɗ��
����|w81@��f���#�'�*m��<��7&���1�����?k%�O,o}PǞ�=���8�'����dJ&2L��g9����<��s��$:dHIP@�/�H:1L�Ic,��X�.�����.�I_!+�&\7��j�O���*i�i!T�]����!�A��B��G0���|�4���&borvp�ZJ_�唐����L��/k��hh�N�셖�֚�@�d}�Ģ��a
Խ���,q[�c��\�o���=n���1R0D�܅J��b
�:�"-�y]�Z��Āܾ>L���1z|S���^��v)h��m�V��Wy�$Mv�����A|��m<������~�
) 7�կ�9��\f�߶��>�[:Jc}���b��Y���܆ u�7�]"�w����ڮb�ްIl�����`!n]m�qBt��q	�N�i	�}�ma��M6�I+@��)ɖ!6~�������H������+����#ҭ�{^�m�>E�O|���>����̟���HY����y@R!=��|=���Q;��}ٖ�"��Z����烈�8O�pB������=���y�E���8�Ħ�hK[(������}����j�\=��Hc�b/
������h���;���,M���.O�~���/]j@줡����x�#5�6��F�ʊ�p"��[����s�<ܙ�"l�J7Ё���-�t� �!q>�0^&�/$�u-nWbD{��
�PM���S�PUU]�����v��N	�6��O�Yê��,L�-)E�uSL))��0?bƔ��\g���O��Ϯ�#���g���u��F�H�u�iݿ���E-���'���u q�}c��=����ut<)Gvh��n���A�����4�����~�~�q"=/<]b�	��Zw�e��m"��?�o�:�fϱ�M������nʅD'8�DAE������&f�%�zE�y����lm��3���v��>X1�fW���ַ�T]�p���k�fqs.�����п��]ϳ����Ta��a,��x�#���RrF���-�����-JO�~*S5J��v�\u��4�>��� ڭ���c#v�PL��L��.�ݾ�%:Y��i�=p�j����W��L����:c�����?pc�m��D�a�kt�٤��:+�!c���mԆ�����_���@gmPHz�"��|ek�\7��C @٫���iź?������.�^�z��נ�b�QcM熮rvSj�U�b��g2�h�Cep��1�% HT�����;����GZ��z8�0z@��<��:�����j!��z��8&��$HQ!�AQP���o-:�p�� y�]AH�����^"��$��m�VCyj�1��{�#[��e�V�٘�i\�)d#0��$�nwݸ�5S�}@`0邟ؘb� ��:�m�\��Y�qU$�����57L�H�ѿ�(��I��%��hÍ���K�)�.�(��W�M�/���o�*l=-h}JԟN�SJϺOҶnPV�T1l�k[���`[�'7�v�g{�˯��~��4P���!#�Z�H�G�o<N6���ΈFY�V�he��T{7n��L[A��K$k�I>��+16M����/(�/Ў�����9�9����p����_F`���l]ӆ<*"y!���u$���A�I��Dq�3k�JI��l�g<'���׈i�p��	4؉��Lǣ�ۛ��iSښ�(��>ޣ�8k;i�Stc����e{c�`%x4��X����Z�����2j����yn�~��y��1nJ�nݢs���k� �^��`�Sg�QR�K�]!\�P
����]}�ck!N��g�z�c�I��;�AF�5&
����(�@
_��T%��9�����-��m4�I�5ed#�z��Z�P�-�9�]ǙI�
l��]��A����Q@֖ȶ�ma�%����N�׿Qo���4�6��V�DYhYk�E������V[M�����4idc달��%�Ѫ|���&������=2�҈��G�6F��~�9y�z��:=&n�Kd�������G�>�/d�!d���(6(��妬u���v�J:��b�^7_wݬd>��<%V��=�N���4�R��p��);
�'�N$�����$B�;���1����c��x����f#��������R�ytB�nPhE�P�@;�$��)Nnκԣ�e=~?Y���Ԏ�ao9nE4�w+9Ir��VX���ǣk��~��ǔ�6��ͱ����ߘrD���b��k3G[DT@F}~#`���v�w������v�~�3��>
�QR���\�d��y���U~�t�W��Atb0S\ʲ�e}yS0* 	����f�v!�Z� %�������9�	��`�Ve��2�V8)|!BF��O�j%x�:?~0�l_D�҆��p`��+l�6 R�D�`8���[��'l���q�Z�FS(-8YlW��� �b��mo4>^AGV�Yl:���z�~�H@K����>�f`���r���D_NK���7ܭ{��[&�][ڵ+�59PV����9t��1���D�K�m3ی���)f}T����Ps(���	��E����UHI�v��C�����iZ�kj/�d��o�� ��Bm���}���ͺ#�Y��K�����5+�H�.;0^��B:��fl�A��+��ڻ+ջ�zCs��}���i�X;L�nۮq�]��?�L���U�H�z�E'Ft�=H��4Y>e�5�_����Z��*��e/�#U���!��r�Ed�1����Z�a��1��Ƈ�r#Z?���0Ɛ�t��,�El�E���Z�Ē�j�q���:�!��E�����D�%,Ē'��;}�Qs��%2�L�3��ύ��y�	k+x,�v�T� �]��)���Zh�X�-�2�+�"A��X��v%�b��BJ)��Ä�+�@��5����Wb����y%�9G6Y����<�U���z3D���6�8'�6.��}?��UC#��E�2����lmry�u�[�M{��)�����rB����F��u!��ϦM=	�?]3�7�~j��s��M��S�U,�X���Ƶ�s�}{�y�P,��VD�[��9;�eh�8'���
�W�ٿR���:������}�(?�鯿�WL���x����P*��͗Ж������Ǜl8�Ūc����<z�ẝ�����j����O=��i������N�)}F���C�k���?a��,�@�rSU�=L��8m{���<���K!j�Y�R"�<<�g:�8'ɲW�A��v��������n�`�Fap�QV���<�e�/ܒ�W�C�Nɴ��F)5��Ug<�eL�:�-_�y��ܬ��I-���E�֚,˸��@)��Hc:k�&E�`�AJ��`�[�qΡ�&�s�,k����²ls<��� o�4���i- ,�-ɤBf9���2����V\��J�"��B.�Ht�bJ=h�l,���E�7���,��S�\c�AnX$Zh�tckm:69J����6��=����j,����ϲ����y��A�p�d��k�\����0��
�h�\|�Zx��S���K�n�ma��U�ke�O������d�u��F
�"�K?�Ӆ2���;�?v�/��gQn+�)���c�'m��^���5��~
H$\4�S�K���������>#���D�y�ߧ��)�-���{_o��D蝟O��6K�޼���>$O�Z���uٴׇf<�����������^��k��M����/`l��
;�_v���-e-�a_Y�>H<5����lj�e��k��y<) -\D�
�;�؆��������*�}�I��~���r6��l�1�<���+*T�Up:
Ȗ>�w������J�O�c�촽���>��چ��m`"�����z=��� �I���Ly��@���&�`�e�|�β*�u�^y!��S��Nbzc�n(o��!�DJ��ƆrԬE)�ڿ�1_�5xE^�rwZUUh�1�4�����^���"�4R��Z�U��$�*Y]�s<�3���@J�+�ʒ%Ji�KP�Fn-�P��>S��(G�؈F��T�� �UW����G��`��l�u- |Kxp]k���]�p>)��>O,��	�i[�L$@�����A�XfTf�3�׋)�8VƢg�t-��AF����Y|-Ѧ?���Q4�T��\�GD������p~�͉�N�y���Ɇ�CJ>���zA�͚ �ۮ{A��$]�}�t�ܯu���]��,������#޸�#�^�~��`�Ǳ����H1�M��U�y�7/y5�6a
J���
�Zc/�O}^S�d�bm�6�yk����$�ǵO�>�T�m
MjAwl�- �~N�TB�k<^���lT@�k7��p���l�qhN����8�?�ƨ��;q�/%|��qwKY��~M���S��C!v��7%����WKf*\-۲D��H��R��ण�e��w�E�^�UBۮ��.�����/������MO�N��gg��QJb�$
e�9��*騖�S`�p��
�E�4��uh�'�{U�\�B�ȳ,�5Z(��Z#�l!D��/�
M�,�ucH��T��+��
k-Ƙ��7����y��o�P��;Aa,�ՊŲ�xqq���V��)Z�,�K��T֒�~E���G���k�n� ވ�<P��,-�d#8Eˇ�^ ���a��d��Ƈ�Uk����߷7�7KE��G[�Z�_k����&��s�]6�skpv8`l���n[�[�%^6�|��]�8U�dt�؂&#��5����c?,�[�?І>��&OT�J�f���;�bgMWa����+P5�m����^�3��wJ��ǥ�AS���}�bՙ������n��=%k��\���GEb;�g"�$��窡�l��>��.�ۍ�U�=ѡ�(ݘ	�eqSD�Z�oo3e�SҷN5A�i���.��\]gq��17@���ob�:��4�V��䥐�2�n���`~��`��<�/%]�`��hJeU�x ��:�w�W4�}^��s�v�e�Ю��KaU�x��u!x_���(}^���X!c����t&�=�B0�2���0Wmu�6)����M�WS��G�1�/�F����(�d2��Z��s���yC��$�n�#׈�7ڪ�(�v�)���<!N#��qgggc(���|8�0Ơ�j������f�FCZ�R���	��^�ڽU{��<�8�7������/X<}�i�cJU/�kJF�$�Zn6�p�zӴ����p�V<��R���%�����Ǜx{�Ns��?�@ek�p��ƨl�D�]l�s�[V�΂��޾A��9Чd@PD"Hd��Q���}{�>�\Uyj\"l�~�ឭk�_D$��z�8�$A��TC��!�J�)�`��K�c9q�Aય�T��[g{�������ХT�(��p�7��FA(��X�E��4��x~u�	{A!m�r��I�����i��*]S ����[�P�)ݞL}eP\M�.�KHN �Kp��!�w��wwX�]�;,.Y`�e����[_���9SS��LO?����T7�����Ί���	��$���L+�z��ʦ~��p�4��7�ؘ2��k�����jb�C�\�,Z���"�ٯz�p�N���b�����]q9����G�Nu�l_8�/8 nYesk���G�i����q�>����%�
]Oy�|�����?�a���\6���8\��n|G�~��5-�0����)��c@���eOq�u���ebEF�|�5[Zo=��!n��q�Vz������5Ze��dop��P����Փ�3�G8-<sT����K�,m����)�֚��˴��}�b���X�u=� �-&vm�4I��M˚���ڼ��ɑIB�]��y��tJ!��FY-ÚoS�b�:<�`�}����������R�MX̼!�H�*��4X}A7BS�Z�n������[��6�z]�Z-����UW֓��E���V���
]S��l&�s�M-d#G��&��	�����揀�>>��s�@��3���ꯜ"�׹�ո�/I]�XtYS}&���{[��(�)I$��٩'��?�@��Ж�Δ��VRB�`ɨ&n���X��)v��;� @%27b	.9�FA6ȵ�^\z�izx����jaw������F�s��E*!�E�������Ƅ�3���Ra�^����u�M���Ʌ��1p9O����L�P��6��̣��
S��:[�1�v�/�ӡ�N��Y���dq�i�钼���im�|	(���R�9��*��Ìjdky��X4&!�q���k�h5�֙hN��%'��p�2�ŷh{y$�#��bG�[��B���O�{��ρ�vRٌ�:�7���i�#��s�^�_�Kj��w�cm�$e�8��/�..�����m�\t�0�d��^��d�N{D~��E$d~�"���L�p'J�"�3���]�!36���[<@.���՛�y2�c�E,�����I�xq���_�r��۬k��HQ��o�P�	�k�����BVŔ>�rPi8z?4% �O҉�G�)et*
J�D{E��g/�S#8���O:6��LwP�H1_��2Z��������n����˔�ze#��5����jd�[��q���G��/Yf�똏��.�#�J4�Sj�.�j2x�ַCN��R�r	mP�� �g�<y��J����==�~�8�U)WPX�PlK#���U].�^��#j��٥W��s����̚��]g4�� ��u�vt^_:(��Ğӗ�%��SBk(�QosnⓁV���eܞI�#��%b��Gxx�΁���L�H��*",�x
�����smf���7�J>�
�����(���=��y����y �n����'��k~�1��/?���9M?cZ4���X� ^�!ȩ)}�����Ȁ�b(E!f�8	 ��������U���}�,BC	-7� ��<�h�z�p`�|�%����dq�Wqq�+5/�5�(��VV��_�bIwK�1�Z{h&L�v�Y�������E�'��]��Z(�����ġz���t��.]ΞV�M���t��r����f&�tV�ۅ�j=y��3Q��"��k�J�����Im}�북��y5��$	O������ �c�;`5��'k!���S�n��R�H�Up�fC�!b0s��:�4f+��fu�k�4��\D	�0G�y��)-�N?����H��
�1���� �F� ��)BO�R$6@v�0��X ��]�"��H�a��?-��q�v��u��]�у��W��z��Gn�y�z~=���%.�0��p>ho��ǯSy�hߙ������aV�sǠ�L�8&�/ߦS�_m���u�p~�|)
w��B�����V�*�����#�5� g���-�&�K!�{1"5�%�x䜷�)�;XX��}�66�2C�&1P�@��=��Q?�ݶ�>��;��K>�ySH��h��0�a�g���Oѣ�5�pW�� $ʉ�2,5S�!?��q������I3�U#^5���
���&���L��gQ�[WzKeF��¯�^ي|#��ɨ�H8��ڈ�;��u�k�ؼ����\�O`���#���"���F�k�� 8�X��5_u>������/�L�<v�\�i�y��B���L;���ú���]�,�+����'vOQ,�/��-MĮl�&�ݯ}&�mY��Y���p%V��=���t_���������v8����9$N�����o"�r�F(����ٰ���c|c�!֊����>,�������i�Js���i9ܴ��Ɯ���!g1�iKu���3�������N5�|�*����-�~��Rբ���ygM2a�۹�P���x�x��f�f�5+.7����T%I7`e�|�t�nk;֗��ǀ�����Z(b�Ob�N�*����,������� q��g5;$��;\-D��T�)
N�l�,����D�%��+j��� ,,��Nڸ��U>+�� ֠o;�g�3'VH�G�"�f�ߌH�&���妎1��dv!r�>�G��6����eX�}	j�_|���UwÍBN%`�n�p�(zv\�D 
b ��Ze���	L�#�**1i�,�b��O�����j3q�[�s٭��B/T�?_���;�,�P9�|�I����b�f��Ȝ��k�X�f���2�r�2<�l8ɧh�SA��^(ͿW�^���|��J%���?aQ��+Em��'�C��Fy�)�	"�g��2lmdO�~���Y��Z�Y����z��V	�J;�63W
.=)���3.�4�j�T�:�o|"SA�`��2B��� 4[���x1i1�u׭&�`W�_��N�A�[�B��47��ANZ�|^�$��-}m|~qv�����`&�UE��l����S@�[�q��G��Q!�z�n��G@��f1鼋��D��X^��^��|ڰ����FJ�%�W&"�Ϫ�$[^��̕��Fߖ4#����w�Q��ޖ��������p7�\x�ʤ���z�,4.�j�sl�������^$@��g@H�ݙvޝ���r��W���^��ϳ��9�og�DA�oab��P�շ�d�qK>#Ě�aqy��!�{�������k馊2�F?�����V���X�<~+3[�����������}����K�D�N�����,���:f�䱓�y�ϯl�~����L(���G*�F�0����$�%�d<8K�^S�.����G��X1><�Z�$��:�T� nyh�2�*o+�)@/�!�`��_���[�]��o+ �c�M��gC;Zں�)z�/U��=y��gQ��x1��諸⋯&]���і��[\��w����= ��.U�����[o���-���������Xo\��m�o��M�H�9���>SwT���!-�����/��82 �^����ϋu����(�x��Z� 5�8�4��e,�F6{CW���Y^-d�ؤ�`��ѦT҃S��O��*/[Vǲ,ۇR7��Gs��R
�F�O�l�����dG��� ��%�8��-~�!5�D
��o����5�0�� �5���F3�CfZ��<�ޑ���x$CQ�kH5Ç���i6s����_s�V�$�����hjPU��2�/���T��ɪ�۴��Q͊<��|>���ACi��H�jiq�ަc�C	K�c$�����t,���"��|t�$���G��u�L�wv;�_���,��!Y�������X�*�v
2��B.�T�-��[ujuGA&�_T�io��ȿV�M1�#
|	ޜl��_�o�'V>2�٩"�C�����,�TC�l��9%��v�~��\�7�j��c�F�= �JuGGǪ��ޕt)4��0;Eg~o�� Tc���F��Y7�a�E�gx�����ȶi/�~ͭe����o�P��=[U踏Tr6�l����(j�Ϥ��c���*��M�Ӛ`C/�:ݾ���d�-3/����=_V��⢾N8�5�[VG�2�f/��N��$�<h�Nh�-I��*�	סџI����Xv�֔�T����T����y�cw-�}y+��l�Q�m���y$8��6�=g�/�I�ᇟ��ͦgY����㇁R�4��:|�	�XeG��O�$�ݱ\����O=S�����M�\�F�����X�M�~�ͱ	g�:}n!%q�_0v�H�[,�N���w���8S	u��e�S�25� ��Y�5[M��:�'JZ�d(�f�B�0��>�&0g��P�y�L(�}NN�R]�#�O�i��R�D󫏙?T+��դ���Tx8���**(��)nY��6w���nb�G� ��ٿ��Ɗ��Z�Y�X)�S�n�VYdrt�yh439�D���Y�l�[(63&@�OCE��b(pu��y�I��ÕJ�S��%D�d5a��*Fq|�;�ygH���E��՜d��߰�)l����q���f��'ȅ~Pۭkd뿋��}!y�-�@�M�XX�@�{�$B��4ﵘ�0��t^�l��wA ��2�{F�D_�I7E�T�&ag����G���3[��7���W��	�Ӵ�
�L����L�)'��;��TV���{!�+Pc�y�n��?Y��+�&�N~6�bOh�o,3g��sL�@H��	j@�|��տ	�m?��&�NNX��=ԝ֜f�p� �$�0�Pg��A����@�?.w�O�0��(���f4^<����}�5b����XW<��Y`�ˎ&4���p򸎙^#	����o��/�q%j�=b��������2
�6��F�.�e�R��5NV��<�-���G}�(�9>�La��T��'��oCj�V�O�E�8��*0~-��������Sa�0��<�m��:�j)7���O�o��hȉ%�a=�n�������vvF��KN�_!e��\_[���D���lBI�ߐJ�Q�
��52�]�7"&�/��WNz���k vwC��0�v>�(:�T�)w!�;��q��X�S�Pu�|�K��4[X�oY�>�Ͽ�u���e�jM�|=?���Q�[a0Qb�̄g�_��{�d\3Te����?�Y^"ѸL��+`��:��؊~��L�O�<�/<�����@��y���}���GgXV$I�X���+NLm���
.��=A��ū!�m$a\$� O^&���y�go=�@'�3�LG�7hg������j�_��[(�Z��Ս)�]Nx�ǟ��<)5�-�Ne$��MK!�J��`��ڳ�/���[�9�8��̗#���o��Lҡ�8L]@s�i�M�~���UO���+����F���C��U(?,\��?��P�/NU	���ǝP`E=�5��aЕ�f�%�hU�;7�+�-�jj��@U��Z��2��Ǆ�����\}�?ʰ��ꀁ�J���x�$���g�=>�\>ϋ˶�G�|�!�Fx��-�I̚!n��=5m�����WOl�
qz�6v��C̦�9ΚX���mU�XfxTy��ЊI羚�ԥ��hF,3�6�1���_���sA^�z�e&��
���;N�z���[o{��h�����$�v��V�����O9��tP�rj¿�v�&����uV�vX\ԏ�Q��A�L�K���[,I6B4狂��{�,{a�,L��6��,����ԭ�"��*(�o?�y�L\�u�6:��Adj��J�Z e�x�<D��$@�@����� ��`2�/�G���U}I���
3�!�!N$��5ѢH�x��1)��"���k���sp��~hxa�m����y-L�IW8)����G3�:ByCCJ�L���������=���k5(��F�dJٔ�(�����Շm���3Bv�H�q��y�����:�b^��Aqr�������(�h�e�ty����V��L��f~]@�Wz�_���A&�����E�>���[�#�(RӢb���~O��d)!�?��Dv�Y[A�v��BF��a�3�_�\�����t��]�Sa'9Z+(Չ׋�k�'��V-J�o�%s��tw���rCJ
��)o������vZ�n�v��O[E�����rr����X�wx�Q�M��'�u�	�Љ��z��	��ђ��2�}\��S� *:�
����i��_�j�t o?�́�D=�W�)ͩ?�6���)r�v~+���J��:8��aC�e%OMse5U=uFV�z�m�iEov���_��D[G<��=}zK��뎷����"�n_�����|�Kd��5ｼ���%���bT�8��<���ɏ�ɯ.�j�g	�:F���$����r4 ���5��\���D�K�1��I�I�Ԭ��Ո>��	P�s��MA9+f{�V��_W=�d'm6E>�a�'����v�/Sq�.��F]�!Mgs�1�^[գ��O���HZ�L�҃�R$�UI)`�5��V�'�����:����O����TRrKnL����,���o)��kUx�;OOx	0W���6�t��Z��贗�A9Y��\��=�����T�)+O��C�Kba��l�9B����Ɨc�?fv�����! �������eW��gu9p^F��o����,h7����5+�g���Ex��O0�X^<�4����EunGid}b�K &�1�Hda���վ��0q���Z�1B��.��u��[��q(��N��6��t!H}���ؚ���|`;�χrDؗ�̏ԧ;_`l]ZE���n<�s�q�t�$M�[֡k���;e.&�8,
�v�0ݖ��8t����NY��fi"�4����CP;����0��Whru";�����[�y"�-���_T�a[��K�������Z�!l;�8�L�G�{^�O"%8��ٓ��B����>+���bsm	c�_�۞+ �M�u��͛��afb>,��)���!��� �r�gx�<5l��5���=�D=]�T�����A�v�}�¦�i�G��}�f͕��S�,v�K��/��H�È���#$r����d���D�� �������^{�9��Btl$$.L7G�;�"g�K��W`�_�����Ri���B�\�8��O�c���,��dM|�ٓ��Ou}�����1V��w
���~�����������"I�{O�����:)���ea�BK\�!T=n^���~7�)ҷ�s��ӳ��mLXO�g��J��U<�x�-V}���t�5��7�s��@,�W:Y1��� '�7��>��GI�gO8�p��cW?&��MN�}��N��ٺ�2�o�0����ܒ�}����}�}ף����4���4�����{m݂� #�4�-?Cb�u���kI�������#��,�CW<'��\/�EW�"�MIf�^���u9�v���-��p�V;z�ɥk��ꊭv7z��
��w���߶�w	m�B0Nk�� �o3�P$j��S�.6'��d��]/ɹv�f+�?MW2��Oq�f�@��j���IB���ǭ��aEkN���YU�M�t�I)�-ֵ�+�q<`�����c��$8+�+�]1�Y��4K�����_Q��m��p�<zS��[��RV7�''{"ޛ�o�������G��;
�R�wƂ�`�M�S�?Ԯ^�6��|��,�ǉ�^������Sb~��tc����R�xc��{T/��?d�&�~VI��F��ϮF�^��U�q�d5�N,���1�_���8���Z���4�kQ�׵1�������j����)����,B��ŉ�e�e&y}���-ÖS�2W/!��!{�?�a��f۽7���W)'|��C*���|E���v=̊�⽳��	��ʘ�݁�w�:P�sh%�.ⶤ'k,�-9�����P�p�Lʐᐗo�g�ؠ�QjǿK�M�s�R)��%�{�"y��BԔ+߼k�Ɩj9�0?�^��Nڛ��������^�#�O�
�_��9U�>�N��]uRk���#���d����%�-��/oA=E�����&��D�C�1+U"qm��(�,�ݪh���Cg�Y<�e�-��	��#)ˀ�Tg��#k�4G�m��u����c2����ǵME�B�4�~�{���4IU�w�]�)Jz����5�k�2����=��"����8�_w�_���v���JA�+S=�\t+�e"�\A����7o&u��� ��$\ؗ��B��6O=lOl	'���'�����GV]����ߜh�i�qѧu���e��3Sٸ6�SM6�h�d�������B��d*�gU�����!�А�rr�Fxz,y0��)1g��� ���֥>�t���9�d�Q�dL�k;�n��F{�����?�<��S'�<�øn�f���U-}F~F�!0��3ڟ�v����=�P-C�WG��uy^ X�$�%b9�4��.�V�3���L�Ե���W������yx�oz�t�E�q����(�g�Uܘ?ԁ��p�?�!�Q��{������|P0���_&\�#��4W�.סWr��&ND��Ŝ���; �a��Ӄ��x���{�����ǩ��'߬c0E��3s�FE���R�R�у�uQ�Oi[^ƹ�ٗ�����֓��k�k��~��=�v+v�"݋���H�_�)����'I/!뙀�|�27ǏNm,I��>Ò��j)5$y(�[��Xˈ
 �����e��$s�+��fQ��J�5�Ā�!�/�%w���v%W�	Kx>�d��<�JgJ��g���Ԁv��4��
B;��,���E���g3}G?�Np@�ހ���ćlg�	Ȯ� ��=�l��N��x!署_��݅�6>��g��t%Py3�o'
bbt8~��[��ԟR?��/G���㒛	w�kR00}�'�,e�ld0����1S��æ�:�WBߜ�l�b���bp�:R� �=<|��J ]Nv]T�hO�"Ãu��*G2��t��|�j�W 	���X�hzif5V���2�i�i���11tb~d����|�0[�O*�=#����Y܄r�x�v�l���w+#$����S5mjL��BK馅`��#��+�����L%A����T�S���Jj�>�����nwl9$MOOgr%Y�IP�-&�-�ɏѤ#���Y��}��]$d�P`�W�ڞX�2���T�Q�6q���]��h�BG�ʴ%�0�0��9�n����}{�=��G�C��z����g��ef��-��h�P_�.+�������"��5>�a�rUڛ�~0�����p��9�3���W�ͳu�˦��E,#�f��x�b�u�G��5�,���rN6L:����.AՀ��.<<��I^��1TW�9˕�؉K3�*%�Z>sr銳j��fU�����$5���f��������X���^��bxX�a�3l��7��n�[¸e(A�\?M������?X���Kl�����rT�z�OX.*-�"	z��wWo�;��k�K���L��~z�"��)R-JX��P�w�zp&�SW-U��v��^���ϓ���ܸޢ�`��9@���7,�&�I�����4���+�V�4�H�e�#Ԡ��m,Ы惫�L�%L��oķ��6���	�����*��FD�NB��_=����<����&ASwo��Nyp�w�7�/#������*^�MC	�MO����􌆢q����l����)�s	��~5� ���3Rql"�i5.��L��O���EC���Ϳ@TØ��G��A�A�)��s>#,��#}[UȔ�Z����02���.���&u�����L4�,�zXM��]a4�?3����,������;x[�ݡ	ƌ������r��ϛNo�P	�݃$'C`�Ѝ�m�x�hNq�a�Pmx��g�>�z��[�xY�ݲ�����W�O�1�eZ�X&
������ƑG5�S5����)5UGv�~�\���'1���	46�g��3=�1v�g�m��E��2Gl�S:@~�'��gO��ih٦�� o�q2n���d'��6%2~�%SF$������$d#.yC)RƋe���sq\=�.:F_h?���z�Z��u�?�Ѝ`�f���H��"QzI=�q:�8
��8g�lŏ\���<�Z�[hkO	-�_�÷�\�;��ҤL�!#oY?\�Λ�����-$��Sjf�����xX�k��n�<�7F3gt���z���Ocmq��8�<��0�A��h�YX�qȋ<��:�)rę
��˴b�h+�[r۲m4�~��'}��w'##��:�ww�mA�S����b1jՏ�1-�ts՗ʠ��~����ĄO��eɊ�r�ᢇ?^*H�U>�@�Jd�s}���he�͜��L�eI���>4�,t����e�s)8�-�'��6�I�oZ�;��Qg�����C=;U�=v������{�#��-q_���%��h��{77�_{^�_oj2�q�Ѿ���%�ى&����R�>rڭ��v�	�	wq��cl�~O�%$��O4`�쨻�����4�u�H�~�뗯� ȳ@d�������C������E.��_����,��ĕx�e��n)�̛�F�1���_x�?�1�TM����6	}x��ϤZ�a+�T��oU��|�*ȀQN����#֐#�����Y�􎠘<p>���vi*��0�(��-^@�j6ւ����O�����'ν`�E�!GEe%�� &@���:�Ѡ��B=����qN,�Z&*�/��ޅfjE����]\�j�4�9��Q�ϴXċA#=c,}���r��70�Ã��&����+䜾��.�~ 0Ao�e����^��p���ܿ<u��2?cF�H^���#��撹Gʌ)����=�� c���Yn�J��$Wz8��eLO;��&Ч�4�M��21�㣱�[���y�S���a�.�qy>�S[�1 ����R�aq�yN\��Ŷ�֎IR��� ����̀�annn>j��u jnV�i��MĴ�/�#&������ϻ窥��L�>�5�(O�kjۧ��o�5�\:b�X���gH�t�
���:� �׻OF���6׿"=�ԴҘ𿥗>��Q_��ied�N�����q?��kg1<��~�:M���}�Lr^Y��qSF ��#X!3y����y��oa5�i�ی��?Q|�cFU����A����:IR��z�ź�3�J�+�e#Y#:2w.��&h��^�<��h!�ZF�"�N+
_�͝\��Ý�:q/CI��P�-�ə1�1�%O�AfT�oD,%��HP5շZ�kY���M����b�����9��y%����	�X�������(����#��х�er��e>�Dq���(�~ҍ<��	/����PP.�"�jջ���>��w�޲7�%���׫/�+Q���mY�~1� ���q������J��2N�U�3�P>���������b����¤yqZ��sݷ*��+�4 S���
�q�l.|�)DՠIޡKG�m�W��2yH��y�����0��q[]����V��3>z�2��yO����=�JM��{=!���Ar<ؕ�Թ%NC)����o�dm����>Bg����'�{��f�-P���8Q�B�b�h�xҽҬTsV?Py��d�δ�MF
ST����zf*��];ټ����Q۰��N:��>,�Ĭ �#�.����K��@�EC9-�ۂu�c�k��Z䀹�y��9����V�Qvn.����5�u�Lz쇰�P����J��|�)������~(�5,s�QΜ	�@��ʳ�R9���244䙰:��9:��9���G������|��Ź�P��:1|�S\��|�&�ظ0�t��w�SQ���h��^�E���4��PXȊ��~����H�7��l7Q�[����Ô���M�/]+t�WI8��9�$� �p<���^��7����:?��a�5l�D5��y����������t65Y�%l��H�l�>�M�5�
��S�WV-�m�#t��++�B0�3�tGҦ��<����،n����0W��6�IMr����8(7��i�P\A7ݠ�K"�O����fE��O\g�|t"��i*yQ�I��d�α �[ӡȞ`�7~�׷��Fi�y�V�������=�+�F3Q�!��~p�Q����O���,�����a��.*�on�1j�0Ó������a���W��ll铥�?.��U,q}�'�m��1Q$h���ab�D���φ���j�I��c�j���}�<~�5�C�z;��@3Ev�.�-�����kgU"�5Oj��{����b,�Ju�k^�ҿ{�Zͺ$��m���~����F��V�Y�k�\d�{���t�%_�Z������;�.�����'w��لGc�k���ۻʞ�=��#c��-�P��b�j:r�eF�2��Mz�""���]�٧a�sd�)��AH6/L�����u���cyE�h��M�rG������7��á���5�i'_Z�y
�cf
}���0�<�JWI�B��c�'����"vNɐ�S'6��= �)}@�����|B�������|d�@'�+�"PS�{y�pa�#��Yo�ֶ��<�
�S���y�o�!�������#WWם��&���va�e}WOO��Te�7: ��Rο`�Ĝ�䆃>���5rH��M���|��H=�1^$�x7H������3h<�-����S-��mHT�gCx�G�$�P�(��hDz�넋�΀@Ŗ7���g����1���ڃ�����#���L*�	V21���?箫U҈��ط��2/��k�h� ��m����6��)�	ʍ��{Z�a�����M&�jGGc�[�,;�q5O>�O�w����q�Q��?�B7���᧖/����x{c�.z�^�(���-ܝ�k�;�W���8��9:�o��\	fNz�:`�����"���O#�ԝ��[��S ��v�6�f��E�<�a�W[�O���(����ia"3VS�D>�������ּ�״;@>$xzNxxxވ'��3�w&���⏀��r��$1�ON�i��c�>��m�>9#�g�/R������a2vC�Y����Lj��(���s�t	�Lh��G�NGW� ~C*R��T��a�+�ġ�o��q]}Mm�Ic�G���^��}��F��<��ý�����/�'��� j҅�E
��9�9���L�&��9'��A�^�w���R�^������sG� �~�ڥ(|�+��t��T�5��JG�|�l�nGx^���j��j�F..Gi��&�iA��t�z�ѭ1��Z�ܥ�є��T�dA�*���%#�0m�j�5)�ue4>�Q��=�L���^�'���d�.~׏SC��?=nc��M���
Kz�>Vq��w��KQ��w�A���È �?�&=�`a�2¸^pIj�����tq��ݨ�a�cJ� �����3z^$d_|{;������g���k�%����	����_Y�,���N/�KXd�r���MOο�6y��ksB��V����^���o�=Y��Z��M�b��|!�aaa P����'Z"�%��ǘ�����-�p񘇸�
'@��}¤˛~@�ِ���QVV�7	�>
O�w�L��_ҟl�}:c�Ed�=����GXCzC�&��/�~�>��\`��<�[�T���c"@Ga�E�A�������+,;�=,�������;%r�&�G��4����Y$ybu�?�_,�1W�M�dD@�)i�E�>?�	����hfH�� �i*{��Ɔ%�nU�,��Q���v+v��~�4�lo�tfύS����I$��T�-s��z���(��F���m�q�i�o����k���>���-�rTIUՖ�6�N�c�T2e^0ϙ�0H�6e�x�{�lf%��9�����rs��-ܧ��� W�Aq�F�E�7�������A��{�<6�1��Bl���>v����~�Y_R�`�����gby�`��B���+�j�us��K)?�R]��r>oV��ng�3y�+��i�����W�ڿ���;�.��v"u\����V�t��:>O��ϱ�����,&��^v�.�3�q��C[KuUM��$r{]<W��:ڻ�֠5�������M��18��Z�>E�&o����<���ޕX�؀e�]Q�G0|��= ��,$�3�I��U'%�~��y�e7m������[�����f���/@/�d����lxl ��uunwf�~g����#4K�a����D�ns���3#��i��������!��:�a�O4�B���S�Gmk��#�M�ph���wq�C�SNƜ$�L3'����jƊaXJĕg��v����l�l�B/�F����B)���~:z�@+��ŉ���� �AO릟0S5��Yey�hYN$�������BԪ9B����
�����("��v��^�!�y����D��O�׶ �{5�M��i�+�w��>.ҷ�`�>�i-�{B����6��TL�4~�K����X�0)���[K<���,G�Yt�G��&��L�I��K%e�q�,j�dI���,��������+O�B�Ef ���=ѝ��x���1�UQe���z#����o��)�^���ĵ�II�����`���|�����9}f���ذvE�b-�^��3kڪ���F���K�5��ӽnqE�:i����+<��2�],���q�	���:�>��~2��C���ܧ���f��6���`�N��M����3��q����)�{g�m��,|FH��j�D��)�����?�v�h��&�7��<�pnT�Zz;�����~���bާ'{#����%���:Xx
D��m�7��4]��?�}�$�!���H���W���t�ƣ�� �۾nd��q�s	Fݠ���=�
R_v���������"^��}gI�6��4��8��j[���k�>mv����]h��`�*�Q���P�j17��ԅ9�m��Q$�PQ��������ll̈���?�y#1�
Y/;�j��-��S幗őF%Mj�:��6Q�:a1Y.QZ)r�������C�}�9�*��s9AP�N�I#�JT�����P��F��y�A.iV�@n'�r����K�ۑ�k�`T*S��^��[J|���	�]��_`^1���	.{zĸs�,�A��)ֺS~�/��ALA�l��;�������On�}��*�C��EU�Qk�J`�<X)n��>��ɦ̳���9�{��s�Ǌ�帵������׫�彈S�Q�k�*H�Np��(���齊7Q&��;�	�!�b���`)#E�=�|47>0a��Q�%�eq�?J�����,������nW)L�	E��[�X�	t2{����Q։iV�77�M�?�0GTƶz����g�NC�������������[�o{�u�<�_4�!Ї�\�k��o,QR�����n=����;q���v�ۍ�7O���5G��s�;�-��	g���"��������է�?P:w]>�<UK��1�8!��;�r65�8��2rs�ZA� <HM[���{k��s(����nm������J/�j��t�d��'L�
T�('�[�p�ooVC2-�1\g����S�t���Q�9��-���͑�
����8U}��m�"�ybJ�)���(F5΁ǁ�#_~Ƽ���,qܣ3U�|lX�ֽ^�Y"���_|�f�N@��H_�S1u���yIώ�/M�(m��sW�����&x@<�z���>��(�4�����j&�2�^�ͦ��kB<���|!��H��?@G�F��y��ۂ�� ~���Oސ2�|@���BTYG�g!Yb֜a#  �p~��W{a��]�zZԣ�m�~����)2�ת�>�$��U��V}v>~��A�G閖'�p]k��k'� �¦^c�����Y}���F�ʀ'R�c��?�f��~2��K.���K��1�L��-q�x:�2{�����K��feǴn���w��;Z��5�&7��\�&�{�1񻌺�h�����D�?�#L����B��s�Ղ.R��^~�+����m&nb^�����m�����U�&
���a�r.޵Q��."w#�����fp�Z�\%d%VV�/k�,8wC�A7rA7JJJ&v }'��
W}�&��7�Ho�f� /�T�>E|�֏鈃�ql�.��R�����`$�=S�'�3�L�lhV�p*�ǫ?;>���l��?�cXG\=C�h{�+O��_��K�����v3��O��__́��w/�ҋ���
�����_C}?m,�f���m��>��`� �@N���<ϑR233���?���������6���#�9���,��7��EAY��a8VS�a�́}4�ߎw�a���Oꦌ�QG�]���z�#����}{��y�fXC�;�*T7�тZ�8L�Y��u�ZW()	�%%e^E�̢,˛�؛���?w�����x�֎w��(�̥��y~��o�c<Y_7Ysw��Ҹ���r��������5�{���#��;���o���?��1J���|A0N�����{)O���˧�T~?���&S�F�I��Q��^]��
�}�5%�����c���~u�>��'���ϣ��{>����)�BA��b*�`��d��YZZz���������}�;eY�RJ�Z��s>/a2�1Û|���e/�z�e!��x�`VU��� ���?��Oy�Wx��9v�ǎ�Z���*UU1===���g<�����������I�0`o�y��XG����/N.����Ez���(h��w�QY�v��~bl�)u��g�A�|���K)����|����ŧ=/�bˡ�<���3�T�Z� �ISj4.v��~^��|^U�M��$��șm^����2�����41��4�F9z�����E�8�'�;9!#r�(�\��UU�t:/���_��<���j]�r�K�Ν��[o���?���$I�333b8ǈ��k���㬵�‌<�у����8F)E�V�Z���?��x����aaa!?���YYY�^�ߴk?�|Vp�J���2)9���$In���8�8�ep��ٽ�G�K%oRC*�Q9!J�N{�`�[ܴ��Y�#���0zףh�������s�G?���nǺ�*/�%��� ��Ш�ǅף]� �Q�~��A�y�+��cd�ey[GdtTU5^�oǒ�yCE�pSH)5��L�+8�g�N�d���
�HӔK�.������_����������5�������3�~aff&B�~�/ʲ�m6�(�u��ߌ�v@&�Q��(=`ss� ���i��^����6��.Ƙq�ըxn2`�����Q���ݰ�	����*T�a:��}!��(�.����[�؞`�h5��qJE8�J��!t�q�ޕ���a��ч|[�`�����iq���@2"V�pk4��`Y�)��=J�
��4I P�pvL�wӝ=jQԽheo�.,JI��>e���7��R�
k,�V�$��QR�#h������t���/G����Q[ȉ�;��� kB
		 Nb��m0�pm}	��x�	�O��%q��,)QR���k�m��w���G�1�����[��������x��h��k]�2�0$�c�0 �"�0$N|��&�h�p�<:�ߣ{��uJX�P��fC�sʲB[����wN�B
1�_c�(���(����'�:�U��9�n���v�M�z���ښ�����~��h<�j�2�<ϣ����9TUE��i�R��n+,>r�?��h�i�5ƌ�nG?w::��M;x#�`��^�x�
>��{<{��~_�����.�1ꀷ�9���Y�v���@"�wj��mS�/���H����IQ�l�:t]��,���*MRT���R�WV��)Z�@��5��f1�$�L����L�\('Z7�(܀.Ӿ/�Q�v�Z%�J���9K��4�h����JS0(r�2���"E�2'��qLUi��4�-��-Z�i��X�Y@"���-+_��m�׃�\��qٍI��
�֢��O7�"������Fk�|@��C��GS��8&Bd  ��wר�Ɣ��4��6�n�7�$�TDR��p*@8�D(�q���@�_��cf�������k҄������'�,���(!��� �Y��3:9)X�\��r�$���a%�Qk�Te��*LY!�D��@
��:333ĵ�0p#�����>]TB�q��8s�;���!n��;�����&� )(����3��H҈l�!�d}{�����~ޙ`�I����;\�J]!�f�F�α�GЅ�@RN@FYƢ�`<�܎�ҙ�7���ܴ>:�3���&
#�*�^�QV�McY�Zŀ�OVft�}�pNH��Z��H���:'���job+CZKi�Z̴���)�$���%JkX'ƛF�ф*�s�Rq��n��Qۀ���a����	���I�b����HO�X���EAUU�j5�UU��v;�ߋ/"��t�q�EE��\���FQ�Q�dm�����d��v����.��ܓ���x|��yy��!7�'ք��;!eUE!YYp��
��IDc�����:~�z�N��dnn�(����N���F���6׮]��s�m.�W}�4enz�4I)�3,H����}p>FƗ�N�pBF����w�q��T�5#4a-��%�[lmn� O?�4��]���l�jL155@�ݦ����v�������_���J�յ5��g���G��Bzv�q��Cb�S4�vm�1�y��
K��hDU�YZZ�����F-��g��'�dvn�Z��l6I��4�Mڽ�W6how���EVW���lӪ79q��Z���-�(Aɐ��scRݜ�9�5�ǅz����cc�	?J�8n`� ��$Q���
���E���8u��_�2G�az��z�Z��u��]�UQ����ҵ+�?��ka���Ǚ��&m���0΍�nX�$���H!V�]��F�я�=	��A��w�]HVe���<H���O}�	Μ9C�ޠ^�1;;G���T�[�l��i�z\�|��W���i��ݤ�m��M�x2[hjq�.K�1$����UN����G���w �<�N�D��� S���N��&�r�=��^��4Z����Qk�QQȠ�ge}Sj�[�|t�/]des�����GIk���h�Pa������(��Y� wƣ��9�v��j�`���q�����v���U��WQפ�����Ⳟ���Q2P��B�cn��[a������%yN�j��S���W^�g����sssT�\w)J�)�fX'��6�Ν������?���K��p�V}�GO���^�K�$�̤�S�,���QL�T$0NЫ��������c|�_���S<��;qH���
oځV���v�]6W��Z���7��?�!��m�s��q�g�������Vx#��N�к���x�w��
�(bym�յ5�Z����
/�+<��i/2???�(E�p%!���"������\8{�7�z�w�x��Ͼ�4��N�!k}�
��"B����7;h*P(n8�����l�2�<#��$EQr�������#|�k�ę����:s�4M���@	�s������=��l�w���x��wy�����t�+�K���rdnc����-�!_>�ډn��Otb��KGG]�j�XZ�εk�0���W_奯���ӧ9|�0����th!��iG(GQ�>R�cii��W.�����Ώ�bee���U:�T���UT�E1zXg��C��y�2Q�:D�
%J��E6d��de�N{���S-~�~�_y��Gs�����Y��F�5�0MK{{�K�.r���ß�kחx��{�NͲp�8A�� P���t� �5�8�MxT�c���[��G�����a���06����_�����/��[a�4M��V�.��n��^�4���N�]MF�$�߫fc����o�s�����O�A۝��T8)�!7Ғ�;�pmy��^��cg��w~��O<��''�C�.�n��(PR��R���i�bK8�>�����˼�曼������o�	�LMM����C�a�ܭ=wG@��at#�U8_�QI�a��m�C���4"���U�;L�N�՗^�_��_�:��;�6yU��&P
E�R+�$	UU255E��!�0|t���?�?������0;3���!�a�7�@�b@=x
��" �݈ �R�T�� �K�b���2�1�~�1����o|���C��Z�BP�Ic|!!H��x�]�D	�ц�������?�Kν� 9y�IR�!��팾��aw=���`9w�E�
��8ͫ���,i6�t�].]�D\���7��7^�ǟz��3(�����qƎ� PX�鬅RD�:��Gg�������_���D-L9�x�4J�m�+�T�$��w����Y2ސ>B��FE!Fk�wvX[[�̙�|����W_��g�Fr<�GF�њ~�Q�Ij1EQ`p�LOS� �������	o��M�y�]V��8<�����Γ@T�%2ӕe9N���>�`�b�8�#º@H�ц �,p�n�KW���R�{�9^�5�~�i�f�|�O�S�zYmJ*��kQyN�^���a�4�?p��~�ÿ������K��'��bzz�@WQ�!#LY�5� �o܏cq/�ueY�(�.����{n!�և�d/F���v���b/dT0J�RJ�<�i�Zk��_��^}�յ�����o����� \�Jk-v���v@��`��: �٩�G������-9���$�E�����J?�s��	~�W�.�}�u=�wߤ�7~F����#G��j����@)_ObEU�)��J���[;��?�.������9u��X�9G����5�~�H(����n����5r*�{�y~���1���eU���Ag��BQ��H��$��+��*�<'��	!�ƷG-��ѹ�/����w��]� �Ա�J�N��\�8�:��6�����~
A %EU��A�����Zgi�ӳ���o�}~�׾���#dU�����L58m���(0�&���� C�F�c"$U��7��[���!kk봚�?~���e9Iy�9����,1֢��w$�e�xqC����4e0�������x������u^|�E�����u�������Z4(��Y_ߢBzY�0��n����������;��H5(8v�8�Z�n��;�a��D�fRzb��TDiJiK��\�x�(�����O��7���S���^���4Rވ��aDE��>B�A\�A����§6�f�lll��[o�?����>8�������i͠C��ќj���������LT����,���Pb�fgg���M?�o��o�w~��F�z�<��E�ք�P�H�T�������n��uY��b����$�N�����1?��?`{c��'OR�j�O�sֻ�v��Ǳ�����c/d/]��?k����79�b+��Guw���O�m���z=fgg�����_��W��������~Ǔ����W�
�Hk��+���6�'E�9Y,s�k=ldң�ݱ�x�s~�E[�5��,q,a(�v�lwv��O�����_���ќ�FcY^Y�o��[_8���0]o��1���U�/�FȀ@y��2/��%I�r��iΜy���M�\�B����x9���;�bx�D��� ��Z`�+�p>�EJ�����di�:A��[����6/���-V�V�t�"�PL7Z$QL,�0Ai�0a�rH+	E���|�#�T5,�?4��{��ʥˬ�����V��a`��Z#ă�gvX�}����Zc�o��������lm�s��	~��.���!a���F���C�9E�B�(���8m��XcQH�U(��%,8k��ӭ'O���f}k��/�9��I��߾
F��)o�wi���X�#D�~�C��D�u���A��׮P�o���ǿ��������HQɀHԢ�I��D��D!$�8!�����%�[[(!9y�$/��Is��UV�VQJ%X��a�|��s����7V�$�؊��u.^���E����=~���S���G����@��$���@E2����TH��@
�#��n�5ӳ3=~���O�e�]�L��C�V'��8��<å�M3�G��_��f)%N��s�Q%!B��K��tɳ�?���������/�!�Y��.E^!�*@ȀP*O��T�Ӗ�
ϔ���r�
K�+��[,^�Y��S�h�\�p���5�0 ��8��E���ݰ���������Z_F"����؆{}o$ܹ_�n�yʲi�������=:���ȭ�����u��Ds��<\8İ��!p�EƵ���˜SO>Ư��?�o���8	W�\�'?�[�~�k_�G�275��,� %"���E�NHE��8�H����� ��K�<��c?v���%Ξ=�����i�"G�������Y�Hց�r�8�²��ᣋg9z���~����~��Ç���p��EV���LS�=J�$Q�p�HF8#1�#�R��l��T���������JYBF1�=��f�s�@�ۥ^o �9�F��z��p}���rL#���A����������o�FQ�|t�#���)Z��Z���T���Jt�	THĠ%�(�QH'�v�* ���Rp���z�Y�g?$�4kujqʠ�'�"_2$	���c��k�x���8PR!h�	� l��YY_!N"~�7��_�>ss�oo����nM!úI��Y\`��@�� c|��@��1q��s輠���`0�^�q����q���]�J���@!�'-H���Hn���7�A��>�e}{���U��8����y��ߤ�Kʢ�ZGU�(�)$��w�K�֚A�K��	��!�9�Գ��u�;;\�z	�����y�E1�ڕ�t��:��FQ��?1~��{����H��,}�J�F8�����9�<�V�ʯ�
��O~�3O>Ne4��)�:�v��( �d��pZ�)B�Z�0�҈P
>|�]z�ӭ"R���h�YY����uB���R�$���'7������f8 ����_����������́�p�p�����-�=<������寿DPK��j,//�'���Ȉ�����Pk�*�d��8�I�g�U�I��~��;�C�P���P�%O<�'N�`}}���ϣ��0�@�N��.�iW����CbP��x�+H��^����5Z�M~���~�w�(M�g��}z[�=t��O�L�8�p����� N�1� A��0��%Rx#�	�Ʋ�iSY�cg��h�������p��,����HqCw'+s�;;,o�����&����c�}�ip�w�}�4�9�x�H��YE #�4�:N;z;R`�48�پ0;Lo���,s�f����O���ԩ3t{]�t]4juҤ��)�7j��P��d�Y�|N1��maA	��,Si������������n�ɳ��G�֑�5�w��(�XG�P��k,΁.*��aڢ��iR#�cvv�Y��`vn�'�}��iΝ����-����@	u+��}; w���ޯsm�����˫K<��c������^x��(p�E1�Z�.Ji�+ʪ�9���0���,�z!���Z���sZ͖�l��t�]Ν?GQ�,9B��r��)���~�]�>���#���	�odhk�褔8�tUp���<�;��~�w~������"Š T��X�ǁ3~c�K��C���1�ɉ�]����qdn�7~�3.\��ԡ9���}��a��ޤ��E��)�E}�mq��`��d����y��w��_��]��?HC}R����mw~����n�R������{�����3%�A��ac�ܽ�cZ�!A��C��fu{��#s���+���˸X$!��ſ���-�޷�͡�9�AI(C�xQ�႙RQ��<�Vep� ���:gq�p=^��l��;o������!̰�2/r_?"|z��?�)�����Ӱ�~�X�	�����\X�������M~����8�|�2W�^���S<}�ib�)������,��%a�C
�42T�A���-B)�P)��k ���dE��o��^h-M�
����I��Ϛ4�A��C8~7;�J]�tY�\��/?ï�����_a��y����������M�R
$�L�.�(')9q�`�F����A�C)I*�0�Ű�!�_ �3��(8q��O����K,]�J-�3U�S�9�Rޡ���k�;>�^#XN���8�#�Z�$�(6w���x�u��?��\�v�0�m���;�)�����S��B�(����y�tn��f*�B��AR���Ii428z�$V8.]�D{����1,�����C�5~v}�Z������	L�
;�����buu���)����/��ـ^�G��D|�����S�B)�
�i�6DaD'(��BXd���<[�m�_�@�&����l���������eP�5��k�;E����N�qt�����z]�aX5$������W�����t�}B��WԢ�WB⌏�FJy�`���A��Ax2�BgR:�T�I���{������$3%I=A[���6�[�4[-�	���h��NӨH_	q��֭x���O�������z���$F�?`b��}�A�(��W�۔������n��pιQ�ȑ#�8 �2{~!�w�|:��(�"�(2zY����3��՗x��g�M�DiF���W7�櫯q��t^�� ���v�����!ay�o!�H�0zd�8:��<�����Hl�ly- �o �o��ҥ�5�
Ѻ`��E�4/|�E��?��Ԧj��M���������q�'O=EHH�Bz[}_;2.l�;�^�A�f7_�$���8��]Z��Y:�>������׿���
y����'%%*��|���5��M���<��Shgy��X]]�䩓�M��F�N#m�\7|Nm��΋�	_���<m��� �(�	�9�WV8~���[��̡Y�]����&y���İz|ޱ��p����5�����g����;w�<�T���PV��j�޺dM���$c �W
�dq~��%V��Pa��_�o��_����UT�n��>!��xr����)X�X'����������_akk��m����KN<3��zL��a����f%��V�P4kM����h�M���ߧ�Pj��S'��_�e��-�{ַ6	���򤵹����2666y�������0?�H{��0*�4a�V^y����Mַ��^oh�pl%p��%_z�9~�_�ܻg��_�Z���,�;���>Acf��KKU������=%	p�������8"w}�G�c����q�;a�f1�	�c4C�Ly�'xꙧXXX��$jNq��s�W���S����ǩ%�a%v�<�A�U�'��k����P��@SJ鋎������SR�ҋ/1;3˵k��)�5�:l	��֚�/;��;�,;�W��
�V�������o��oP"��G*�`�(�4�!E�wD�I �12���B�����누�^��ajj���y�(�����j�bX���w������&Q���׿ʋ/�HE\�v����pd�(�8z���2���YD �g+	���@�AeK!P��e�SNUH�D��w(�g�z�'�x��,X�\����Us7�z?.����������fna�o|�,,,���F�����Ѫ7��@�w���S�D�Sc+*]��R�$�X��e��.1;;˗_x���y���1�`�RU�M�������l����<���7�����Ή·�A�}7��?9�[�!STx��n�O���駟�j�[o�E�ץ�h���O�ԓO�!���y����?~F�̣�I�v{� P����>�s�$������Dy:�(��a�U�
��k���ِ��)���P��N����
Ó�����6��p��e�[���c<�ԓ����~oHM�����~�z)8���������^3��bПk8�ʲ�+�8�9C�ߥ���&�;Ac�A�F4�:�N�w~�sR󵗿J��N�(�0��*}�(�j��49&R��y�a��F;�� CkOu:
ߞ>s���<�hΟ?��N��ZC�� �(M�Nw���y�/q��ӨH����ˬ.�p��1fpVxv��s7�A)|���n�x�[XwCi\���>���2����*/���?�$�~����DY�X[���-��:�/�ҷ�R���|�2
���c�Y���;+p�FQ������-�W����q��9B!�N��W��1/��3������N����C����vE�� dsg�RW|�[�����^����:�F�$J�5`��mj��pDo�C�Xy3�8�v>��*C=�s��a��;l������E^}���llmS�7T��+EF�C*EQ�Q�����-��_�U)��(�i)�Gϻ��N(�;�Xhm0F�� g,�4�8z��C���C�A����f��_y�CsS���zK�e�������n���_�ŗ^��ad$Q��	��j��kѣ�y"�*��8�s�(L��@�(��\�0���<����ϝ'R!i�0??Oc�š�yj�[��cuv!�׏��3=��/r��
#�T�Z1Z��y��Q��ȸi��v��ʙ۝������}���᤽spw�~�3�n�ڊ~��� EX�0�RV�p,_�N�-x����iL��%q� eH<Ԣ�,6T@E��*���ԑ�,�b@���)����0��!/��"'N�@W[[�>R���_��>e���Sb��!	�͝M���Y���ԧR�~>���?`vv����2��"Fp&�굺O_��4�qƎ���ᩫj"�F"�$�cB����&�^�'N��+� ����E�&燏3�v����Cq�W��m�4��W^���!��������H���X��!��THE�!���k��m@ر#|��/�9��T���&3��N�n�ǫ_}�㏝��%EUbF������w0:����F�N@�?`u}��ó���o�K+K��Ѩ5D���#��Ǝ��)�X��|�++J���x$���X����V���C���ꥋ�\�F��r��S4�u�67�2τ5�Nt��o;<�pN`�cu}�����7����?�Ǒ�D*@%�4%C]��X9"�
H��@޹���5��>��e�t>E�j�Ն'�@H�}�!����f9th������ȰVc�=��B��5�(%���E��W�;DI�)�M��.G"�BH��C%%C�# ��_g����7�Y�-$�R�°8��ӧc���v��C�lwv�5�S�4�"����xgo�S/��p��o��a�sw�(k�~k4vf2b?4�F�p7R����nsnq��޷ȣ�|� �n�4S3-Z�3Xi=�ުS�%�����q��q�p����yg!�qU���`��ʣ�ٱ�7O Jz����8}�4O?�4����W���+�a1���-�X᙮��S��}o�'N�ު�2��k�k\�|�C��h���}����m���Jʪ�Q�01�I%� m4�����fB�SVXkX__祗^�����{=:��C��nf.qH%(����&ӳ3<���0��v�*�
�כH�hk�>�*P2PC��9��^�v]Gb�nX�y�}�)+LU�JjH!Y[[%��y��gQ�bsg��,�iG�����5kt������K_��E���lln7�"�(�[�(⬴w�GN���Q�Rb��;�Pj�h+)���f�E�elm���3gNq��q,���n]T�TIc���0��;��V�׿�DI���ׇSU�R�H<���f�5��F���eEY���X�1S^9��Xc�}�Z;vff�fI�V�~���Z���c�I�uvv����R8�r�qQ�%��R�ZS�s�=˩S�Ǝ�d���X�Nk��0�'�J#�FJ�t����"��2��Z��!Q��0�9y�$y�ǥ��	IRK��4%��(�2���nf8登��;��?|����}��8������%m�4�hi!�JÃ���V�4I������R�Rk
m)�y���>'\{�� ��׳Ǝ�U}$�b�AH��?`j�ɫ��Jsz��N����۟�A�k?n��c0�S�����h@��aWVV�����@��r���FlepƢ��*��dJ�WF�Έ�sV��UXm@��1��unn��{�ם���~c��TU��Ld�G�5D���*676��j4��aj��L�[c��ѮB[M�@�pNڑb�+�[3L�3����8&�bz�>�9���?�@��R�Ø�'�Z��u����~������ƒ�)
�.4�2>�c��m��c'Dk�&�0QQ8~��`��ȇ�1�sXo�:K��D�W
��hL5x�K�Qo6�j�Ƶo�!�0C�9dE����9r�N
J]!�X�@T����s�1~C�MڌҔ�kc������;��眼���i���es}�~?���daa���&��-�M�����\�i��a�S�<C����F���j���p��k�"�%"�� ��IJX���D	��F��FP9����h�($��kױ�3�Y��:Q��sY�T�
�q*-�E�_�>��b٣���ހ�b�(
�$D�J8a���/je�T��ǎy���m�FSYC^�?ʲ$PqǱ/*ޅ����;v\tUQ�>��Ӳ��,��3����� �#�H�~�\J��l��de���,�3-���f�,�mw����Qo��D� ��dy��،��2�i7~��<Ash����h�CV,�Ҙ�����i�y�P����#R!A��t��NPk� 9���� ��+���iƑg�w�ʜ�*�u�S>�E�!����C;��s���l������u9���O<A*���u�^���!��(����C9y�~9����JP��1C�X1��v�v���N��9�CU�pȘ%�u4�y-�$�4�\�����Ѭ�84;���&�A�V�ɱ��8r�Ɣd�`\g��izXϢ�$��NV�gDQ��SǑ�c��Nc��Si쐄�(�����]�3�$S�R!IR'BO�<$k�*MQdTeI�W�I�I�9r�(EQ����6�0���jr��qZ�Ue���}�V8|=��4;�-���y��'�����\���
c�����¨^," Q1� ���H���eF�5��t�RWTƒ�%Z;$H������j��
K��iJ���Y#7Z�q?���j`��;=�s�v���]�D��NJ�&w؂��<j�ͷ{ir��0��d��^�؝�vysw��~\o2m�ac�k|����`��Sa�#���A���"��*g�%Y�K������q%("4()PA�E��`�^cr������PA@�8먴�ӷ�T�"J#���&/2ja��#�z���`��3ߓN"샷��ڵ�)?�zHڈh4j��9�3�8�^�c�!	#���8O=
�14j5��_��c�TI�2��a��B�6a���V#��(BPT%SSMJ��س��x�(��m_���r��xK�Ŕ��p~����p��q�8���Y�YG(EFLכ�;}��HIO5+��D��ᐾ�8�PA@�8'��A�!bȺ�eU���A����g$�^���Po6���J�����S���+�������`an���^Q1n/�{3�M���ڊ8�y�'+(˒<�=�<�5Og����R8j�:�CJ�0�Q2@Yւ��<xQY��OѪ*T`�E8A2ܡ��¢�#�-B	��lv���7�p@��g��'O��R�0����ӭ����=�bO�ύ�'��&U�z�6�fĳ_~�(h)�&�[RW5�
|=Ш�)H�D(E5�� ��a�/�$*RÈ�A*�ikU�����N���S�i��u�s�9B�0�P�px��^��
�b�s���>�1�%r�}Ԉ �Y��^�3(�����Y�8fmu�٩�Й
��Z>�k~aJa�0�8����c0�AH�P�ٰp^w)Db�� ף�,�#�e��bfn�n5��̥IB^�H	���T��)�Q����u7?�p;��/2�=�i����v��Rjlk��xz�0b�m������������h�����3a�^SzQ0!|-��!�a͆��`��"�����r�Gj�Uu#eh��)B��
�w��$%�Qė��'N'��}׾�b[76D����a�����E���+az�Jy"Pʧ0Ӊ��:�z�&'9|��p�("��R���km�l?"�bl� )MI/�Ґ_}	����"�;���=BI�$$����B:�EI�^��X�0"	#��Q���(rQU�Wb�U�cy���9��
��"�Jᤠ�*���uE�ɓ'y�'|$m��	!�<��'���Ω߿�����ܰ.)Tq�oJ�DQD���`B��X��,���'e�.�J��y�B(F�I'I�����I��,�Ȋ=2L�$�E�I�7����׆��;y��f��G�$ID�UC�R�y)�xX���AK�@JBI538�֣���-�8FN�C��!i���A�)��GФ砫�j>��Y���92���v��Z�P�c'OľF&�"�a5��qk5�������
T�.}�ַ���R�z��;��0�0"�z�.Z�C�'c+�ZL�m���T�� ���E@���<S�MF?&��poQ��v�|͆OqЅf��'
UF��E�X�"��AP�!�0�B��ДRy
�(B*�5�JWlw�>�j��Y��ZC0\X{�a(��_d~~��.��9���P�E	�u�٥F:Zk��Â{E����v�S�ȟ
�5t�$�<χm I�:b��]�����;XEQ�W%y�cmE����1k|RVfd&#�E��ejj�8���3�5n�,}���a����)�$��J:��n��J�������HP���$P�8NQ�_�Ԇi)9�z:�0�	��C�XMi
��t����7�;���0����`WR�s��(�C���y4���`ks��-���AD ���F�]UUA@�$�aD���J{�z�N�ߧ����F�p7܎�uQ�����looS�P�B���0Q4,澵V��c�iOP�%�F�fs
�t:�~��#�Q!Q��F
OTE���CE��U�1�ħ�y�4a�R��A+�������I
�ǵ3EU�1�BYx��(�n���(�p��r+�h4R��&��CY�8��+)����z60�)m�Z^���m�T��C6Ȩ���%yUR���t��"�%�h:�.UU�ɐ,��HK!)���Q�'C1�� ��{q@_�(|~����ǃcl��0�0֒�Fy�N ����ho�TM�^I$$(��`��l)�]օ�Efgf��{�W�󜵵5��hg���H��9G=����.��djf�0�<�{8����5F#C�R�SHG*��IL��eeu��ј�N�R�������+ա�l������Z����������z�F�/�6�;"BI:�6��X8~��(H5�-���QU��43��r��r�F�����#�i�P�K� F(�sƧ�L]$iÇ����ְ��M�ݦ�4�
�V��c�����063�e���:SsӴ��(*
ȫ]U>r"�O�{@C[H1Ե�,AY�Qi��8���ʪdcm��t�<��.��pC�|���$Q�����0ӊ�z=����v�A����4�y���`�l���I8� EV�>gI��~4� ~�.%IJE�J��t�3�T�h��&���(���	�Fs��\����q�T�ѵ����6�憲�Lr��%�� JB��^�0�Ɇz�*]=��+k=]p���`X�\���&	C�$"$i���~qΑg~�V�QO��A�$��\_�R�T���[��f|$�BJ��`}{�n�K+���������_��� r��7��wɅs�yz��������?jE7���k�٫���\�n�?���ю���}F�!��C����PV%i��4�."��Ǐ 3�D� �By��4I<�ː2Vw9k�:y�#�����8q�0��|�t#��7��	K�Kz��as�l0 d�)o�0C-�����M��e�q�~�c�5�ѣ�9��T�0;?K#��4�M��E��xA/g�h676)��f�>��Ȳ!SSSԚ5���UY2(|Z�6�N�K��r��e�vEGüs������1=�I�ODQD��5Y6�9������t�]j�:S3)�tĳ1q�%1�,C(ƔΛ[�!)KC�ʢ�#
��|�P�cC�?��,��K�Հ��+����C ����E���($�r�����ʔ� :C2�a�����I��e�Z�Bk���Yo��FiW�Bd�;;;��]��i� �!�iwp�p�ؑ��KY�X�;d��� c��m-�8��A@?Pj_�o��Eo4���~Xk	I���B���B�X��)�����2]p�M�m�����Vz��^m�j۶m�v�v��UW������d&3yg��>�$�_��*-��Ϊ}S��9
��F��u����[�Km�w�;ծ�PӴQ�3�� ��XZ�ۅ �X1K�S�o�Vm�"H%8Ol�@�'k�-�V5��B��#|�����Ҙ���!(c'O�f��;q���)'9`"9�f�K�'�q����m��4t
�%߽�c؅���$h=� �[����;���ʴ���P�?r5\I"w�wl�(Y�>)�*�Ry׽t�en�t�x��{��◀G+�IP��@>u���	�"M�vD:�ɏ�P^K<��꧇��DELh/H������NG�SM��Q�Vr�C���H'�I!��0�YZ�db�Fk&���(�/u�Y�C�%�aMQ�8%�̞PWV�YA<o�ј%>�T!\=��fE��"0ӈ�����ьbS��I��@)�&ZZ�Qt/h��S����X�t�7<�J�(!/��|A�"��K�5�(HX���a��Ks
pJ���y�����+���g� nj��Ukْq8�bu."�AQ���<1��a�ޛ/1xF̐���^������?o��=G
6>9�N��u
*���ą|��vş~}}8���Zt��Ǟ�PϠ�@�X~�J��;��ϥ[�Q� ��),~T��&���O������m�m]���3H����MO�<LTROr(r)&�©�Ն�g6�~ڵ�μ-�P�*�v^#�u�����:���*s�Ӣ�Y��gA΃k�3���������,�(&�{<t��Q���VB�t?j��T�ɕ�^�E9m����~�I6��f���󮭆�=�Z�������IoF=��#T�����#�+�<@=�+Ӷ�}��ω�ߜ���V�e�ճn?����a��^��� VQr�)oQXEu���N�,|�
(�Q}��i���&���~=QYò�����ӧ���� ���].Uy�m��Wަ�j����9zD��欒��у&��N�SPJ�G�r��I���6-۾�
h���o��_<��c�TfU=#a�3@M8�����6�r��U*����o�J	�eΰf������㌕l'�/|���U�ww��E %+E�r[�h!�"1zV��ի$3����2�-�Bh���jPH��\0�ɻO<���v>��j��� �@`��:���H�ݲ�ÃQ�@)� �մ�v�7�sh�|6\"��O�Q�}Gx��������e�89-�-�9p��Ilʺ=��y�Q�?�T�{����V�/6u���{�ryhTw��KENT5��+���K�q�6β��R�袑	�-�*��m��$�ZN*FA� Q��H6�?6
�� ��Qhji��^/��\p�N,e���qP,`��G���"�UU�Z�����Ӗ���㍐Ab�"����0�l��z
����Ru;RZ˼=�r�gԡ8��M^�ܢ0r�M�=zH���5bU�O]Ħx�� u�7�qV��pB�	�| 9y��;�-� P�N�n�(��Tct��qhp��Rc��βm��eY�#E��$�_�����U�,hxS|���.����@x�ٵ�8�<�uT)=ccn]���U43��u�}]ScK�
T@��klJ��tl7>�;�	d�����؃��Z�B��+PMck�bN ��`�"{��2Y�7��[��X������iy����H�B���5�*J@�~0�?�<s܉pْa�/H���bY��Q����GƋ���G�����v�\��Jp�R7.�1�������9�J5� -�8���^����r-�z$z֨���O3��w�W2�ji������C���0����1�Z��!$�a�|�c���s�(�&��zKv�0��}�Hۊ0�z��޵&hc�EA�֖��;�)9�U���-��Y:k�W��#!i�.�i�f�20��ftO��s�)����g�y>s�}�bB�w���e3s��G(�-��U��KGt�.����R'�z��sM�)��]����@���kͶ券�Њ�x92�����]i��#��F�I�cI��Du�| ��������<�0�m�=�]�-Rֲ���<ؙHp��{Mʐ+���"�����%73�( �ؓ�^ 4�ݔl��d�a'8����� f��R�Q"$��ڶv�%]�[�gY�F����5�E0b�oT�m,F�����'$uF�N�-�C������Q���x�݈���bo�T��<9-:2~!n�|�����Xo_�.�<��߂H��z��F��A>�W*��p�]b��[�`s�a��i���	9 ����:Ic��Uw����!S���u�f�y9�������F���%���\��եɍ�Ό+�B#�T=�铇aS�ᅚ�pj7.���rh���mmއH��RY�_�%���%x ���t/��Z*(\1�9�g����1Rݺ��''o��Sghq`�S]23T妲Z�r�djj?��u���si5�T��8�g�$P'g�,l��m[{�L`TZ��L��N⢗r��f^����I��ݏ��)�����*^����ڮ�����D�2�Y{�6�z�����̾��1$J�!j�n��.�!E��s��I�è�'H'���BP��R�v�7�ٻp�>z�w ��xp�Or��?�����Q� �nV6�^��3͑��;/M�{32�Fߐ��iIMX��;Z�Y>�m]�Z.E��_�瑽i��u
�ӱ(т՘*){�կ[��K�a��_�P-
�)eV��.���_N��{���k
r�-ӿ%'�������c��leY�7a3P|0���Kz�)��$B��hV���;Zj^�v����9��6[�!��4��{���V[H%#}	{�R�$�0��,TS!bY�I(���Ũ�����!���RT֑��9������^U�yź����
�z��4	�b�
R��/���W~����;J;��{b��*��D4�h�T������Z[�lUd*Z�h����O�
�
A�Ar.@��ř��)&��m�t[Z���3��If\y�N�~�ջ�f�x���3� K����``�sk���b��͏���@�"kk��WPQ�ɼ�g���o��-�Ks�ː���\�A|���KTa�	�$�|�\x��k�Ҳ�r�兪@֩�m���U�����%B8�G��ⴽ��|�p<�\��	
��%�9�^odS�PT������K���Գ�p0}c(/B}J��H��w��KI�99$h�S��@�Z(�[_�u�G!ur�jF1č�%�BEa����F�.Q��HR5�)@*=u5{�|������S��&Hz�޷�|٭Sͥ��ɪ��%�@k�Oo�s������ �Z4W6#�ۇ���y��ml�Q�b`Pä)`�����0���"�ǐ��嚻��\D� �Z3k>%����sBMIDL�"�������:w$��2N0�)��`gS1���/ф����Zd ��V��� I�"�]�V����ыȇ^�t`h�E�3�a��%�7��q�̫p�E3<?����X(W>ޮ)A�cjo�ֻ�I����y�,]z�}7q��nq�v*nq�l#��^CÈ��n��?
�%� F7��������R߬�WP�NQ����"�*��aZAL�y2�yY�"�:�8]���,@
�d�Nj]S�j�]�>y�����5.�x�Im%ٷ:�����W�:fmh�c-����r9Id�I�RƝ���㜱��a������F���xS�`�)��X��%�=?�ז��-�@&2�f&7��Bc��n�߄6���3<��l5=qgV)���{O -�=�<��r�xW�({��S���$�u��"����7��}�i��Y�s�1��_�[��>��h��q	��;ق�����4:QW<}XxG����G���AQ=�����nC���M�G���Ic��o]���g��y�t��e�MphI��y�dgP�Hs(9��Iʡkr�	���K=�f҉��]Q�52e�s���o�*B%d���l�[	qV�K,�'���Np	<4Tא��)�4M�BZ�ٖ���y"��y�QsZ�;WS�+���i�6����"R;XO	�PgĤV���i]��_�_����O���Z���׾Q�ב����{0'%�7��/&"~J�	mԕ�U��Q+��E?�ƀ2�����3aW�n�|GofEf��D$�l��7>���7Օ��V�X;���J�}�?��H(��_���`J�:��K	�� ��
�$�ɻ��xHϴz2>�A�7N?D<�ÉfqA�j`ɿa�#� i-n,<WK�����~V��`�������RBß������b�mu���tIh�%���e~���1f�P�pʺT�2/�og
聼��� �mZ+����|�%�$4g���E �8M�ut��t�3��[���ȕ1W�u3<���_����j�7%�'�^�,v+�i����e��0�
�&,ZjM�f��uO�����[Li42��5Z��7�v�;���2G��H�N#p��OA�\��G.�Y/���J��If 
~����"n�࿩��2;ܷ�����V�J�3�04�D�b`����;��vK��ګ�m�XR�/�ȥA�
�*�%T�@��1u���ޘ�U�b�r��^l.���#ɴ�l﬌֌	|�(����Eh��Ÿr'׶??O%�Ӗ���%V�.������.�(�,C_�r���J�����v�����<W��WZF�f�#`�QK��a@F]������B�߂��R��f�9J�Fb1Y�ɡ���) !IaO�G�:lP%�"lG��TĨ���(�S�-���o���ק�o��6���3!M��[�fݚ��i����|�钸a�*
�'f���h>]��e�.��Ld"��/����e4���ʈ�R:��Ҫa�L*a�����v��;OQ�����w=��2}�ދ�3�C�����\�g������ڟ��V`٢��a�H���U���;J\%EE	j�t	�LW>KSC�"�Y�b���Λ����c�����J�:� ��*Tm(�;2���0Vq���A>���9�G��,'G�Z�!�AW�U��|��?g�{K&�Vmή�� C�3g��[G�A#�G�\�_�����|�W�bӧ	��Ԝ{�\�i-�B2�����;~6�6,O=9�YF,ܐ�J
�EO��i����r���(D-��M����L���$�J���D��@����0A��=��l�gu�(��E#�ώ���ʄEE--�dB���-�y<�S2�#��p��hL�Io���`_� J&Q2Xſ!%��W���Lڌ����R0"�wݪy������w���F��m���Ÿck�LU-���)���*������O�;���e��6σ��o7~�W�5�~�^;/�"��򉒲�#c��k�I���]b_PǷZ��vf����6���-P��C'|�w�V,��)��||���l\�L%,s)�HJ�	�v��Ĝ��ʫhL)�R�����ʁ~c<�ĬIL{Tƾc�c�`J���z����()�J�ޟ�v�D�)����s��-�{Zg�?��x?���(NN'Z�[����'�j���A|�o0+���et����1��{G�6Q��F�lJŚ4,L|r&�XTS`��F�智Bǁ�Q�sx,\x�d�m)��~�������*��Ǧ�w�*"���5V��Vܜ��ߨ�i;c����:Ҹ���~�.�磡��2�k2\j0?��M�[8�T��I�E0Xr]�(��V����q^�ŰWޤr`���pN���)	ɀ��X��nD��EC��̋ȁ��d�c�Y|�A�{���L�l�⎜�j�Qkz>�O��k�=d�i�|}�ñ��!�h������w���z0�'�NR�q
0�ᒎz�OZ�YНz��A';�A�9�q�)Y)w�|��˼}�]��c媈�&R�A���f(�ŔJ�D�{;���v@u}�}��>. �6�4)�-�w�T���X|�miۢ��uj�)�o�h�53��*J7'�-î��)\��+x�J����a�0�g�� �:���[�Y���]<5{��wL)
E�|Y"nVB����D�h�±�g�+�[�+C�ɄEZ��崌�,s�o��k��_�[��c���Wi߉�o��l\g�'���ۦmv�<�Ƴ��$�S�( ��������l�3��=]3��~>��\_z]��O�L����~+����I%LĦ��(�*e_F؁+�O0����{�r\��8�Z�kp4MP,�A�v��e���bx&��i�NP�y���W(#��U����.rh�yU���J��J9aD��t��$hKh����i��f��������c��������2d������$��
N�/f�|R)xS��}����+��Vǽ�iȵ���� ɻ�Y$�kW�8`�`�[~Ϋ��:��Ϡ��ddd��~���s������J���Q�r��v(�U�4N/��,$�\���+��Q�1�����m�G��O�W�G���q������#���|#����+��Y^�;@��	)�r�Wx��`D�D#��\�g��-�6gfd�;"�ܹ��뗶��I
R�b:���J"V1bb|{.9����%zg{?��A�y-�i{�7/2��o��l&^� K/��P���^˶֖s1{n�b��xU9:ϊ�7����"����Qbxu`�050W	/��t�lwȟV2.[��qo�l��R�Q�YR# ����h�2�/���^�?.Y?��M������;����?:³�!����Ef���
V����j�����л���6q��n�֦�8¦������#��D�v�?yd���9b����˖��ng�P��;�c 59�tW����RN<S�ٔ���ŧ���c�q�v����v�0c��HHK*��;rckw���	�&�;'�&�y�|��+%g@����#��⑻,�H���A����'���-'pr���;1�{��Z[�Μ+_E�
IL���`�K�`������T���q�~�k�ٺ����>Z���Z��Hs��������������p�Ip�)��U[��������MrI�.y�!=��;;�Oz_�v����~�����h~]I���Mu>7�Ϧ�l�)#��	nOPmG*��zp�*z�xr��nW�����/aÍ@��2��~`~2�D�!{��E���T���ҙo���w],�/��OJ9�}C`�6�~�~�n�cw֞hl�%�ȹ�>6���N��ӂ7���{��x�87WW4nBԂ��+<^GQ4��Y�Q��K?�>mi�
�N�y31r�A6Jȍ-��P���o@!��*�����:vvQ�CG�ٗ_w�+��E��V�%ӧ�B+��|n��z_�D�^,��~��������֢�����co�<�˷���>��W�NZ�����9%G�)cKU�RX//��^�a�S2Φa|�ʢojZ�v�(�my<�����/��QlS0��|�qɳ�� �x"�{�����BU��w��r�L@*���)B����u�;��Y	��q���B����c u$�fSSS g�t�,y�$00i.�>�KQ�7�dYc�g���	�GL���u&EYG��[Jcj�Ec�����&|v�s�W������Q�7˫��{TQ�}�����ka[kW��<���n���g�-&�*�)�*\�?{<\�D��-O������"g�YË1���	��_HI�Jl��f���á�.9AX�[�#���m���i`t�f#���d�@hvb�!L�t���o�g�b��U}C�B����j�:q+��N��R�Eb���-�W�yR�"�]G�=)��a#Y�O��?s��ZB,��n��4�����3�j-�����:�R67q	x�ē(S	���3�9zZ��QύEGk�$���0v���ZY�5���J*��C?��;�^��R٩�˯�u1�����L5
��G�%��쿃�R�g��`7�����\��n�zL���p:�
Z&b�h�c֜�c�������F4���D�v6X�ЖT�N���땗��o?���f��+�\!,�r����w���m"�W�S��!%;��[��,��,Z	�8Z�.��c/�~�E�q_��=^��tp)��ږ�_v���8��}|лx5" &�dN�8�y�������	�K.��`qq��\FȻb�(�gdKD&˥���~�����?h��z�W�U�P������j���!��_-�Fս�D�x�ٲO��f^�"]���n�Z��	����;���"�/"�e~7������������=}.h��@BEa`b|*�Z~qOo���B��;�"������HK	M,���阒��8�fm]CK���L�����:S�(�%5����9��֚�C��ϑ���s���/%�]$�N�A���qm;�i��?^��h#��X̿J�L8�-�qo�^Ϋ[��Y,���5z$ktL�+��x�,�p��u����x��
�H'I45-%����$�z^���&N���<�JXo~��7eOj�ַtHyU�<�T}cd2СĈ�􉤋d+1���i�U����ϝW���5�\3���>�5�OS^`��jq��H��9��}��%k��ӹζ߱���S\�Hs��&1���J�@��e�3�?>����qd���/�DLcMmk�����H��B����02:
�A$@���;w��f[�eT��H�C�@ѯ�N7/,/%dF�e��Y;�ye��wlǛ�p?��d�"�^��/��G�qĚa5Ͷ�i���U�F�$���r��:.�ő��{�=��Լt��bn���ez��/�Vj��t�\5st��Sfq�q�ԯ7���l1���`��P�|I�~�������E���V�~F�E�&����%�2��i7��s��K��if���2=��5�@��r9��m'�^'F6&�?38����N
Z, D(�+m��<*��u�qAL.sdR�jjj�*'.Y��=D��HD'} �����2���)-�����q53��w�^�޻>������tkRQ��&�9�%{�n�i�i�q�$���'_���^׼���&��&_��z�����B�R���#��9p����Ϯ���+r����ͦ��΍G������~�^���E�0�+C~�<�(J����XE۟�xT�����#��Ǐ]�����1Ŝ�K��p�5bH�g��w�hr������qu�x�߯����YrR�YXQۏP%��J�H\W������%4R-k�HJ���d��XX8�oo�����OU�i���xVWu:�w^�;�ř$ry�x�FvW��:)�f�\P\c��\��I�\��t�w�C���7�J�1Ɗ�F?���t���:��͏��,���0�pp{��K4\y�課�ې��ǘ� l��#��L��1$��h�5v;��6v?��v�S�*�4��w>�Z�a�2����m��\��3R{�<���+���ﾷu@Ƿg���ϱ���_qdI?Y��[d�l0�y&�����2���Qa ��G��X�Y�S8B#1>�#�ь��A��l�Y�[�}����q�`��s�NMa�����Xj0u�D>g7�W�j~� -I`H�1+(��Y���q��w�t�̊+����s��s�*��ff15w
&=�/�	��V-��1�a�dbR��H� h)�zo��6�kN~c|�F��Ʀ��Mc�c��r{��q���#�ѭ���qE�r*kú�)�S�T���@	z�8}�yk�h���m��@U�٤�{:~��
���n_L\~�ˊ1+ �GF��彐lʻ`D�6,LL��>N�>[�ؓTn�h�˛}�e!���l�s�����`���t�A&�Vho�_6�Օ�tҶB�$\Hq�b�PN�ܺ��N��0�SK�f:�?޳>�>����}mnn2�|�b�kV��ye�A�H�aj�?���5����˓Ҷ��A��m9B�%#�ӺDRRM24�B�����5�|�_zf��yD���&r��$��`-ffr97&*")Y��gL� U%^a��Y�"_����=��;����&������	6���im��s��t\M^ٍ*U*8����1_4�fz��w̤/��>ٕ��>pR�M��������1g���
�L�1~��)�5~�y�EDt������z�O�H���Ԧ�ըX.;EfV�l<G��^�(�娵c�V��WM��djz�i�~q���E�����2M�����OF�I�i�$9�M�+�Q+���N�s���ۻv��	[�%J�� �k�Q'��5���Sl���m�,>_�t���MdxX�W]憒+�(��[��Q��n��Mm
j����bI#���l�N�r��WM|�񎉧O����td�ʩ�f+��uHA����
ɋO�[;#!։6�{#l�jv��[��V,'�'
n�F��5��+"�M;V����F�(&h�L?�|"-XM�LY�x}���d�=�*���\5c*B���qL��]E��xof��J�ԟ�h ?.�"�7}�%>N����]Ԛ3\����^��張"'��L��܊'�|߹��0�+��O���99������G������ʌ���57��-�� E'u�^N��!�%�(��̆�� �^Q�p��"����?W��x^���K�h�%�Յ�3���-.2��X;��~� ����&ޝ����A��W2���
{eXl�.޶&���Ɖ�?)	?�&r�[I��MN������;;y��8nAԅorL��hXˤ��~r/;DF��oЪ�������j�W���;�B\�K�o��k y8��jL��,�#�"���\x�Ig늛�G΃�C���گ�Ǆ�)�Yu�"�ks�����鎮y�r��_>��D�L�`R)�r���!�DL|��;/���*�h{8���7��fT�"�G�(mg�c
$k���@��!�!�M�?�����EHF���K�:�h*:�����jQ�U�=��������ǭ��!��'fR�u=������x#qNF�w�u�w��%ʲ�l�W|a祵�k��_�'�lҙM���a#$��?��ou��my��a{;��]v�᣹�wt��1��!@S��(0��ȵ�H""�q��V����b�^v�"rhY:™�G	)q�0�|�<�ZY�
13�u3�E�UMB=� ^�؛5���1�6�ö}���o�7_vY/�׬��<���@@ �ǟ���lll���/�C��s}�=�}^�4E!f�^aǓH3��Q�őgC�zC]��3Xi"&qArI0�n^9��+���5�=������������y��4y��<D�:B�
�-!�㡏-.pſ�١�c�{<�ؿ-vYb�&A�^鏪�^.�Z=��+.��:��GޯB��ƋYZ#DPs��pi����m��v��j
+&3���ӎ��#**v�%&����60�/�b=�9��8��JFrI��Y��m�3"焻�� �o\|��`ؽ.ц�4��"�������sI0�z����e�~�����qgW�Ad�C�|��t�
}����N���7[_C���4�kk�V~�)D��4A��.*�xI�-�����#S�=�"w�������z���<î���ѕP+5i�l}{�n����N~|�y	�Q���y�*;�$k~��J�U�=:���T�ՅQG�f��H���d�
��=�U)#L���b��
6N�6��%����޺�x;��vzb�|��e�H;n��ß�o�6+fs�(_���O���{0O�~ �M���l}ζu�Ox�wt�j��a�~C�\U	2�4� @�H���/����P� �z{y\���s�ȆqXG%�
^�Q�<ߟX1�,Hf׿����!W�q=��3�QpV��Ῡ���C���I�TVt1��r��h_��0�W�@�M.Z=-��â	 �1ط]Ĥ��'c$��<��������ו�݂��nK\���rv)-�b!Q�ҡ���n����7�7h�aq��/Ҋ�������>LF&�C��7��p��Ӭ�PF����!
.UT̄ʤD3����d߷/���EX��$�2��y��%G��&����Cf��=W�Z'x`"���~��Q��j�[X�$�Z�6\M�J��K���O������f�%��=��-�~F��D!CE$86�MG2<A��$w�V�����l��cHb`T`�Be�&H��VVy����[AQHb�;��#��U+��/���X�8�LY�'����?B��,��/��GRɖ`����I�d4P��c� d������Θ�_>�{[�_�����D]B�>6.�|�����̲E�RԚm0R/ya���	d�,7S4B�_�"vr3�2�a3�@KV�|7/?!�}��Q����4�w̢�Y's��RGb����.t3J��:��v�~=3����v��P[��n��:�#�J��~��K��Ռ3��7)D+Iİ��d��B���nGiu[$����/]��q��6������W=�	A(��y�e�L3�A��C���~9�����Q��Hz�w6fea)��c��*�+~x�혁�6�5*P0�WG*B ��9�q�Eo)�#�������2hj���l��l���na�W���������_����BТ��m���Lh����US�ne�ߛ|�:��ɚ����uL� �cl�#)�tDk�a/	��"]i[�׵3vq�����/2
��E�!?9�=LM����&�-H�� �	{	;!q�{�Rְ�?`��͆�F�5��4�w>����a:�z���8LQ5�!b�!�� x�/��=1++ݮк6���zi<{���_b����w��Q�7�y�I����E�У��8�{�%���]�+�y|�*K�9kG}�	$�����9�Q21̦!4/����p������,+<�s �!C+Q�H��*;՛ښ�=b��db22*$�����B����y
���=���y�S�S����m���l�w�/=����43fmp��mޗ����iD�r�qT�g�?c����m�g�C�/\0��黉�k�govy��WFCV����,$��z�Ⱦ��("�|�PBTďB��]`�խ?���*l��a�Bd�/+NF�&"��Ѡ]
�G��ɣC^iow��ư���E(x��/4��3������WF�V��]SK+,ΰ�߲s|Pe�����V��U0Ƭ���u70�t<�;n�X5Ե%�"��=RN�Âo4ng�e��`������c#vc�g�D����5��Ad���C)�����{��A�0�ߗ���!P$�h�W���~�9�S����'����"��x��<'�*]�fϨ�Q��C��bޤc�2���I�p:yGgG��yK#���uF�U�<0�xA
Њ1yp.��r���J�dL�-��p��1�eä�ˊ�
��!��_��I$�{?�S=U#	&.��$���!�_�b�K�9���W�@�9�.щ�˛S��dVkܨ���'BX���D@Q��� .I.%<a������}C��8Ȕ ID�H�uG%����V��H�8t���C�j��� j�|5�0L������#�,
l���3�DREG�AV��F�����;i��^'�����5����yX'A�K�P���D$ �E���S�TD��KbQ�D�LOZz*�o$z���%k�� ��Q�s5����iy�{��J�IY�FGW�r3a�8�ZH!š�'�B3E� �'��y��"a��ı�#�4�`w �Uo�,��3�4D��'�ȟ:�bFՑd�"p �u�}�gH��Ͻ_�?������^l F^J��P�.\���V?��/6f�/l_V�  Wb�\�N�,�Lfה�V���3��G�s��'8٪M�r��k�C#qM�0`���ó1�9E,������@x�>t�XF���D�"X�B�Q��a��A��������%e�O���Qp5C�b����],�9�@ e"a�cJQ�G��#�x�Ȫ���@V�_��8��G���owD�v��  ͪ�K�&h��+�����iR��;��`q a��M`!�`��C�}ioݲ�֢H�y#Ź+�	�@`ׄ��Ј7��a%���/ز*b�?
DJ�'�!�`k$k�������-$΀X)��(,�g�+��ua�]�a�QecW]ݼ�o���ƭYH7��W89Q6��� ���+F���)t��Q����q�2�j
W�z�]�xC\~"�`uڼ(��b�D���bF�8 ���� �vT�E�(��]CO<
QR��E"9iC��v�.�Q!>dE.'a[]k��̰�?���PFV����M<v����hSe�E�+Ⱦ��x�o��w: &������@����Δ���'m_�J%���Ӆ�S'q$!c��K1'��a�-�--�E5A�ej�cJ�J״wktޑ��(������R�}������/�����̟mc�����_���5�`}�g}רZ�\�osI�	Ѧ6&����JqD[��ǋ#.ki��"GA���H�؜l��`�������(J$�6l�N&�-�e��Z/�(1]ɜ�y�?��q�{b9De6�`���\�p���@J���	zQ�r������ Ѡ8U;M["T��ڟ�P�`c�0�8cS�5lk�TИ��aTa���%��D��2�Đ�����!J+��^�(���K���#�d�ŸP�Us�1S7`���Q�Q���'cI���8���p�h��|���
���P�h�'���0��M��ԇ��Z�V�
Y�ߺn��n�{b�Y塨g�iN�`�� @��3n#������HL����c";�A��D!�-ވq����F}�f~�]ĉ��=��Ķ���o��l�h@���2�H� W�V+���rtT�s�������\�N��)�fם��"� �OqD�#���~cd=K����/���IMդ I�k-p��h���L8?�~ڐ��=����&��ɗ�\�6�y�9�2�޻�����i`��QZ�������d�+��CJ��)���~��߫�UÏ�cᇎ��o�Z���}y|�u���Xd
�Zþ�S������ϫ��zz^r6�� ��o��~|
ɂM��0�H�L�iy��4'�dM��V
&./���MG��9����LHP<ʌC.[��ذ���/�؟v;�B�Z�Ӭ�,���9[�=0�Q����-7�3�Km2Բ��ayl������*H�1��'��B�[�;�s2.qT�e(�@�O����u6���O����(�h�u���%��<�j�1��7	����F���'7sO���lE�N1⟥�^k�ѕL��={��O��4O���A��>��l�6F��Y�EZ�i��/�g���K�3|TysL;u���t��[r��I~4K6��[�
nލ��E�Eۄ|^���Q
�]�&��ڳo}aer`<�����f�KL�@єi���wA E��;��c;�D�i�� �X���-�Q�T���F���уKUWR�C���L��m�0�_[gm��J��X�������^���C���������!�x��v�@A���/���Ǘ��<���OQb�SSjy�����s��Jsus{��t����
蓿l��7&/l���G�N<4V�/J�Y!Z7_\�i:�w�9�i#�����VA��b��\�8���A8cFP�&؈Oߑ�5��TXZB���=�Y�_�Q+E�@$�I�X���Y�<w#���EB��:�E=ˣa��)ZC	�ygP)���S�t��qU�+������P9["�-i�i[��Ɩ��RZ~Փ�k]�xUOn0)�����33�8�8��l9lRvt����g���CA��)"BA����P�h�
R	K:'o."X~��tu��6;�����'�����:11	#kHD2�� *'���� ͫK�*cl<"�ۢ4������go���>�>��X��X:�Y��(˩�#Õ��[�S'�|F8��s��zi}�:�9��u�{p��<�����t�0g�*�
�/��B1Ś�sR�XU�7���?di���ŏ� ŋ��d�É���%����7��g�:/���[}�8	�?JO����Eӟͤ��>���C@^ ЅT�	���怣�1m�v�n"@�]ƯQ?Mgv�^Hox8���`�	��c$w��؍�j0�jIA�+zr+���?�2=hiT5V_���h�j�{�I �� �T�(-�*U@$i�� �TiBR��Ti����BM ��""M�@bH���������ٻ�������h7�L��sk����n��lǯ�y?բX@,�J$�Aadx�݃��(pp?#Ѻ4:�9Ws�h��Ġ�4����<��@Ev/Qǩ=�(;(W]��3�gXGی%��o~�a_ |����h�{b�@���%�`f���䀊���i�����03v����/���#�1KwO�uG�Wuu�,�W�qo�G5!�	b�����3�gL힖�OS��0�bes��E �~.�
�f�V����R:���/5�j=�	����`:'�S���G�!ceZ��X��Iƻ�属�W����A��S��ж�O�,Ջ�Sl~d�J�w�<�1�N��)�.�����쵛��o,��cc�zb%b!8e���x!�*��0)>���Åd�ܟ(��"~����3iPg����2ʏ
�ߤ�
��h�5#"��E�F:y���K��}�_=U:�2h���
)˾6Dgp�����K먝y�x�F���$��P(��ִ�R���>A?K�l�Ub���{� jU����]���;a���.��A��"���x'p@������H!'��w����}��^b��W�[3�$���on�otO����|�����g/4���$��ty��q�:�r\����qMixɓ����qM4�1T��L79�J���6ڪv�|%���l�i乂�h�$�eX��"���8����I�!���r#�c.f�޷���P��́Zӽn�d���FxE���J1�Vɲ���xa�� vr�y��}��6N�}o����XN�M�9C��5Ԕ�/����]�T�M,��[�����u]ӷ�~���%����;0��9\n�*R��#c:M��F7����H�p����ٌ���NgY���c�)��4]�}��]w
�m<u{ѹ�1����tT��;/*v8�h�oz���/���l+��g���P�'-����*)V>t�#���$N�/�CG,�Dğ��U2��f��s|���d��k����v����%�I�}?�Z_@%4�,�p�B�Գ{<�{�l�B��$��D����f���?dT*����s��%o���L�1S��_���R��d1�'is�:���$�l��}����H�@�韋��#,mU"�2��G�B��jЏ�d�.���b����&zyo�R/���q�� ,�>�����PJ��7�-��A`����N�^9���V{��|ɫ�36oZ$�;G����h|ak�vp��C'}�_�|��E���#�_?����s��!4דJX��_\�q�)���\�8S�@0�f�4;�U.9R���!�t�j���N�����b���3�Iw˻z���B����<�Q�y�����t��M '�m�e �-�~q�T�U3	mA97-¯���rP��U[>Q�?68�yܨ*���t@(\�����A�t㲔����/Տ�2����E���%&}�s��þ�%����z����$�:x���V�8��&�@�"ᩩ3�7���
�!s�%��Î�&��;BNA�C�/��{�q�������2Vj�[.]<���*_��J��x�D�jm���N�A˞֔���A,����F��v�p�G1([�T J�����#o�=�p�{d������q��NSਚ�!F<�6�3V�b�3o���4#׸2���p�L[�CB�uo)�C1#nҭ�ÂO��G?��p����f�}��~����l�@�O6��)����7Xx��zW�/�ϭ����*��p�Q��xY}��г���Re�r�-�p�/V�Y��+\������\���SE,�4��J�8����ʦ�m�Qmƃ�J>)�MJ��ZC~�]k�*�������x���(0��d�*��W�f��.�Obd]2k�;a��V��r�8�PrK���~��r�`i�A��~gy�� ��d��*V>�bv����@s�l���J;w�I��f����h?�ɿ��L �=P�k���,�a%�J��q/�����p��eU(k��O_�ๆ�E�J�k��C}nKTJHs��T��L�T<K@rK�^��B*� &�}�`���}�L��Œy�-Վd,��82/9E0ޑ�ęmm&����g	o�9Ȯ�se:�m��䟩_ҕ�K~���2k��|�8���w�2����& L���/����l��I��1����/�ڗ�<�oz'-�Gl�Ù��h�'������Q���g�oC��Wr>Ȉx.�ٯD׆�^#{]r҉���%[�&�/[x�:�m���ky����g���Up]�H��ny	�A�Cy6K�.�l�?��|����!s&�~:���~����xC��\*�7e�����Az��c�V7������2H�3б��S����c���C�BY���Dׇ��8y/�lKC�=f�[}k�.^;��z���2'vB��_��I*��BkM��Xw������U�A�������J.��ƾ��m%��M�|�����(y<f���̿adM�k=zl��'Β�`'�9&�o���CC��˲��mr�g �6P^Ђ�L��1�q3�i�I��O�II�A��Y��+T������'ؘ^�H4��?9�+�궓+G�ЀA|�������͙ț�b�=ny�YR��>��>݄`���bқ�r~YQƲ��߮�BNOd�]bȜi����4�S�6�{$Ho�5���g+���JT}�IDl�!y�i�o�
�����A�����?L1�@��w��Q)�e��.�go�(����4M~��:]��j�1 �'x �4N��&.kg2bw������|��|�]�g���tq`,?��dY㵒��˃o��r�1ϝ`�˴|1H�lz��֜I�����(՜
,��b��o����p�Lhϑ�Yo'��	�-2�.�ڗ}]�_><|8��<N�\l� mG7g %G�C78YD]��ʨi6��x��m�I�3;Vs�F#όf���x��]�d��P��UYҲ@P0U�s�>���C:(mx����"u�&��sPs��x�6ڼ������L�'J��p�irf�M+U1��7�����ky�T'�]_��$bfk���#x���O�Z�1(�F�.*�%{��n�!h�U*J������<�[|�S���L}�V�#,'t���GKU�9��67���3`ɶZ�d��/8\X<Y�Q�a&�u��w�����0�|�2ECSS
>�r� �<A��JW����C�Z�ě�S��UY��eЭ�,�h��;e�x�������}� �'��I��ٱ��c��8�	3Z�����%��\# 0?@�t��?>L�^������-�.\�p/S,U�f�	��'�J���4�"����5��#���B��c��ɰ�,��g��.ID4AX�&���8N^<ԫ�ٺ��p��es@ ��0����E�0أ� *aii����������յ��.�D�qZ����q�(���K�ɞy��2��a\M�{0g:fs(r=�H��V��:�?��Ƒ�p���{I*v�>G�i�)�������c�^����E8e���k��8ik�yaq1F<my=N�sRI%���i�c(��D��X��f�[�~�W(]�� \�62?<�\_�ެ��V�m����S����qS-ى�6����3%lR��Q?)AJ.����*$�ǝ�[r�m��`Ri���Bu~d�!�+ճ�gd��_�,��Eإ痌��m*����������GΑa�TG�_N3;��������;��S�g���:.~����������!�P��bxo��eoC&��N�^ʶ���_A�[�wKin�����SQ�8�� 7X<SL�{����}&�d�4�M]�Y��55���w<�2t��@W�a�d$HOH�L��V�<��߁�@�Ͱ��K(Y}D�&ɪ.��n��-�^���JE��b��򲠝�r�펜��@P�F!�cJ�R�P�<}�v�n�,�t\�!�R�W�_��~��߃�������t�ZZ�^y����GCV���]���0��-����v��<vs����,qF�c|�P��%O��,n�*��2��N��}#r��2Ґ�=q���bZ.h�cZ��*0|��T���xnp3��n�hN>��Ͱ�}\g*5u��h��~κ�����D=��=p|��k@kD��]�r�DH����<��mڠ�`$ݻ���\�?(T��,lu0g��6�����e�?M���"Yǌ��x�H�T���ZKW��8ϴ�]�������E���z�4��zzZZ!��cZIe����	M���S����~!�:��.t�DΝ�;��M�"S�`�h?K,o�4���5����{�yLAb�`�j����ԉd��U��=fa���Û�G~��3�;:T�o���»H�
g5��;[�gK���A˘���K��h�7p�$8�Y��������H:�W)��1�����v>ս���a���Ԡ����3o�[�N&�F�Ǳ�8�5]�����=lg��	��/�j�^:���ڧ��y���X��	gl(�;��G|S�͸٬i���><?��	�T����GNv	�z�0��5�(�h ���m�'�9�ZӢZ�^U��8��r���Be]�t_l�&"�G����Aܵ�:���v��h�JX�{�t��ٸ�^��:0žyDk��Z��f�Mk߇}:������~�{�f�3p�W��ά=Vч�-��W1a��p��Pf�ݫ�a���~�b��҉*4��}���^�Ҏ���:���������y��#o�W���cOp�Li?��`�:u=%���A�F��t���dee�/��nm�������`X���bq\�����:�S���$���u�9a܎+�A�0��9�68�Q�M�|@X돖���WY����w�!�,�sh?y	4�]�����U�	!�?6�
�P��V��Vo�D{�M��:����,��m�}�Y��J(��u���3�v`z],0eF�P�]��=����8���^���PdEGGG�������2V�����zMk�+���4Sy����z��͓!M�PR�a��)��s'�?����k�5wH��
VQ�(;�+�k0{���������q��'�gW�EY���҂
��Tpڀ��"��̹����O;�rZ�&�1�'J�}r@R$N_2��WD� ��1�L��M����o�w;��vDfH��wm?ǭf��K�d��e9���4��.��f�!�1�"�1�9�%`��A)z��Z��ʹ�X�_�5b ���/+��]�]2��fjF8�9��ƌ�O��R�0��5y9$)�T�~��(��g^e#�
��מMi�w�Ҡ�,��
��IS8J��q-|c~E]�<==}iT3zQa�����c��H�T�>���8;&�k z�a�_�F������D���km��Ԃ��4|�=O����ɧ�d� h��D�d��:���z���N렁nr΁\�&� >Y�����y�!�T�����NXw�����Pܲ9N7�}Z�G������B�����2gr��tr�O���ٗ ������ �'p�4��	xy��Bh�|����w�޺�L�R�Qؕ����mӤ(�hS��4�O�t�k\�t��;h?�y���0Gh{Q�ɡ�_,/@��!��+��~�EƵR7)����)��V?i�Q�	�TB�z���\�#���w;@�k���	ήg[�_������[OO|"���l����u@�e5{{�7��@Ų��i(r�A=��[�ڦ���J��1k�I!W�F?���XCǎU �� (�y��uv��M9L) k�[L�K�#
=�Ef)��Ѽ�H-�mU'E�]}����Sg��Ʌ.���\E��͚
��;	��OT��ڀ�޷`��%&�ҰRUQ����H$�yq@���[
�I�hU�w�_���6�9��%�H��[�NZ��@@�6K��@�k��=Sɀ�T��譃�_S{�^��:�gj��E������u�5M3Pr%\raz���k���e�yE��{ʗ1`'����}���P%��ʰf�=�2��慠�=>&T7�J��v��Y�ں�zX|ES�_��5kH��g+@���U�ϲ�^f��`���WNK�����-��8�r*\�5~"E��ǦvH^f����Dj�;l������B���}B�y�k�~t�	\To"���8�@�e��|���>R����+����]�MH�_1T���m�6�>)X�t�_94���k�K����
�+]̍��R�@�?Q�����r%{�B�F,��?U�%�q����}��ejm �A��¿>��3�n�c9.+���Myr���=���S�Rq�V�f������U11m��Z?G�e����U�˜4��ʨ��Aғ�2Cm������n��RH���t�v��G�[#	��i'_ļ'���I�/W��``��S�F���-�d���`s�М���e��·�������Լ�n#�	W�_ �+�������{"M��y_�[� z_a�-�����G9L4Բ/N�W[���z��s�6_n���xz��b����[�4a���2�M�bhz���%�� PK   W��X�@M��  2�  /   images/54862705-cc12-4a41-9ef2-e24c01e25159.png�y8�o�7|[�H�"di����Ki��-ɾe�)E�%d/bb�%����c�Qvb�c�����<���{�<|GG�q���������u^t����� A�ʵ+���h��w�'<L��{��q� =%���׊� (gP��%M��߽�����I�f�rͨ�����6G�0.��3��g_P8v��l�����+��8���O�':�ٳL#��/Kc_��\�U���wu~�4�@{\�{c�
��=j<]����˯�U;vj܃H�d�k��ghe���,�UJ������/84��!���Ϳ�˂���xiSSӊUL�G�����4q��w�ou4����7�:V���So������!u�ݻa�^�n��I�Oed��A���h�5�P`��[uG6������7بݠя�Ү����d�2��W~mcy��ˣ�a}�%DE����"+���G�'vmu�<Ƞ!���O:�G�'r����P[�<f��ׁ�'����Ms�V��iE0�?G��!��|�P7O&+]�:���h�K|DC�.��Z�,#z|{��#���u�E�O��Ĵ�H��WU�+����n�/Xo�pgC�J�8K$���b��m��
Y61X��e�_�ɫM���J�����S�>\؄=�~�޽ӏG���͉��D�t"!񕄮,+��E���h?�����"�w�ޚ�x�#�b�H��h�u ����u�K,�%��c�4�_Uuכ��Hӌ,o�f���:�T�[�����b�1~�G�/�ǟ>}b�7�e�w�Q�j�F�wO�x�ެ�_����u��d}�gL)�,XPY�R�K���<�h�)O�-��c����S$j��pHV�0'��"��}d�m��n6M���^�N�v�poi�c��m���\���Ϻ��u���Kh�{�\Y��B�����֥�~�q������K�y{���l9׶�?~|ȥ����(��얰�����}b�}����X<<��zm卑��;ʉj���S�I�@�3,X,���̳{I��O�un���Ȫ�EG�<'XK΅��Tr��j��f�}���6T3l�\��I}k��~Z@y��.����;S�PM}@;߯� �lH�IvBؖV,���1x�y�FR��ԁ�t�A<~x���.k`�̱��l�P�]k���+S��e��ꎿ�?�Bl3%a���/����=�H�i��O,H��V��z`����%�� `��`�%>V�ANZ���i�51��.=4Uvv�::E����?FXS���ZX����99] Z�OI�=w�-��}y�����ə��Hq���bȡ�<Y��>�U���*<��q�Ϯ9���o5aެ����8�@�x]�K+ 	��%#�`����iy��y�B�o��R���'�X�y��d���$���v�Tݛ?ћ��=�xps��g���ʐ�w�1�\Q�呣w*H��j��g��d\���9���t7�����J�/���{���L�G[��bL���3��27��x�v�}G룆�\�/p���Ő1������ N�#���f� ���Y#�$� �˒t�S�s��LX:���,�(�5��OHl�c�u��;��������GF�y��G;�]��x�bf�}�bځ����g%Lnn��s��ߨH<�@p<��%^���΀������^�~L��v�U���y566�M�	����G���qX�� P�j'�9�v��6�W���Ivy%��,7����aڟK�l��X�(H�Y*��L��1�S���CP�8D<}�`��|k����A+ڴ���T��Փ�6Ω�b��>�Lק�����V�K{�̐����RܫнHc��K]]�xtJ��;�,���4p���#K�+�����W�O��|1k=Ǚ(�Z+�f�x��)))�XHĆ�a�w���t�^s񈏒J[����0Jl���\��{+�\��Y�[A�+��8Ų�J6ES�j`sK�ðڗ/_L����v�`��OgɊ�c�i�s����[���ߘ�##�����RZ�X�����c����������Ą4�~���2�{qq�E
6YYJL��Hl��`L�pp���w�ڦ�J��ϱ8�SM�5^ͮ�G٣�.��u��0�X(����ٴ>��:�Y��)���EH�����>k3uh�UYx�a��I*^�=����(š��������ރ�>>>�
��Պg�E�Y� .ZI�N��\B�}�p'ҿVMIb���j�]�!��9+ǵcb!K~y0��b���:��o���fQ�nn7펲�\�e��c�l������������3a�+���s�%e�9,j�ֱD{{�'{��5Үē$���<K�#�;�eH�vwrr��_�Ԕ�⯽.�F5eU�(���H=v����e�Lo%���k�����/8�<�%�����[�s8�WR^m#���R4T��&u�	�����xx�
OW.Wlt���'o���󣛾k��}�n����>�m�Ԑ�4�&�k	�Hi��*2�_���1I�s��D:�L�N6�Yc���5VRW8���Ȫ�������N�sl^ ��Fc&������z�q���g��	��4nw�$���sMiU2:��z8)��$��D���;����y�Z�zlr��mps1��
j�Y���#���4�Y۾.e�{D詁�I�Z���H��GH�������ĢJ�e~�)��c-����)��7攔F..F�� ���$�Of_7=_5�,� �ߢ�r��iI�W/�������n �R_/^�7������o�8���<�.���RF��W>	�>�x�=�(_����E��O��M�pMs��/s����N��0�1�vDBJ*�._�5/�|���ي/�U�I^��HkOsKKCM͕��{��{O��/w*$nR��d�ͦ	���A�n"���t�$��>OTߺ�5'�[�lI����&b[L�F�A�<�ҧO����K����%�ɱ z6[��8�y�Q�V��`�f1raK4ɏJ�8�DwQ����Uz_�Dvk�Dh�.s�Hd��|^�Hx����(��!*��/_:����GP�ٷ��b[���!B6�E!&''�E]�v��}� ��I�DD�ڎ�S��?FGGp�t�te>nС�q� ?�8g�&�k4c��p��#��F,��EN��;=HW�>q��������K�����Q���Z�X��]�e;ƌ�y�z6��y��Zx1	L�)��j�>�����ז8�npkgV��	,�m���Z����I�"`�TD2!6=@�A(��v�n��ZZ�O^p"�\U\�P���@��[}��[\�|¨��e�u���=3�Т��XZ?�0�����[e�f�ܮ5�,�y{��ي �Vvs`����k:&ff;��F I�����LD������?~�uf�b���?��֦]�����w�`������Z�N�S�V�v��y�wA�Ǒ� W}o��H�L�PA�Qcc�<V�|�`,�}��y?]�b(
�W����N�مL���略E��ظV���n` ��Պ��5e��;�Ji�s��4Q������������O�����B<:�+Hao����@���hg���z�d����A�#�@�N]	��� �.�9�<t,���(��I��F������A�Lٙ���#��n��x�~G������/��s056���r>��2�;d��K�SE����s��CYIR�S�wOq�YAv�j��ާ^��D�4�)rs�Y���L���R�i�o�ؘ�lB���VK�*���(5�;,gb�v����$���떺�H�}n�{gL�v�Jp��PR��!g�O2s����` .}��!؄�4S��i��*X�!�=s_�=��W���� >����ֺt��_K�%��h���~�5\Ʒ=�ЀΩ��l��脄ȴ��9�!��3tVx�~q���;���C�Fک���{������ i�cɝՂDjȡ+(�5�]i � g"��K���nF�>Ȭ���Xk^tČ�8'Ѿ{c�c��ĜhF�`��7	w�ݿI�{.�"�R����A`ҶAG����8��g���&���5I%;V2���[�291��S���ɬ/��Zeڷ����kڕ�8�E��)�J!�H���zʫ�|�`�m/��U&���[������La��U�օ�>�i��8Aߞ�<�(�l�׋��I���BCB�So��B�Q�&I~�7��}Z���1�Pj?V�p��V�* {���`�n:�c"��s��n=����&1��~Z23�[6,L�X@���JFFF� *H��V���@#/^�x�3�(�<F��9sR�gy���p�O3�s�hR0l��Ҥ����뢓���]~�ctf0�xק�555��V�c/��N�홲�&2� +��g�{x�<��s)�v5�U��^�{o[���ii.���V��i� �q7��"�AU��t�A��� [�G!	���'�z߿�l$~}�2����?{�[{V�W!���I�(�"�� /���<��d�������V�}�����t�~2ٍ������ܜ_|��w%���{��D�(�K|ͦ���4m#��ͪG��|��C�B~���Ƞ�=u���)xy�N�u�Kf��p����f�V��oF$U�G
�(hj��BV�Y�W.Vԁ�l�#S���&cC��Q��oe8�x��*�������y��I###��El��	�勥7��׎�w��S�`bb����8�Է�\��l��"�Z�	����ݓ_�|@Hu���j�(~�~z��I��)|~��@�q�~�MzUr�>�-;TG	J�=��o�&��$%
�#W�����7sss�b�]���݁�� ���fJ*6`j``��t�i!�R�M%����]�yy�l"�������nڧ��m&~�њ���Z��-�����-4�Ikv�����;(�����z�(3U��6���A�@Dn�3/K5���߹���Ձ��\9S+,���	C�,�=ǽ�}�r�Vtpy$1lJ �EA�*!ː�W��,5$R���S���z�
�[F��������z�x֓�FTގ��$/e��^�w�����̒qA���&F~��`�iy�gs��5�l5��M����.�R��C�I�	la��(dD�[uݗ?�{�J�+�)��ӯ���Ӗq�
ٿ"�����ˣc�y��5$�����ﳂOl���;�7��K��]���Z��L���S�����ח�F�EC�m�f���C
���񊊊SO\k?���p,a�n��W����p}��{�+(��Ⱦ�r}��!�rm��I�]�!e\;�4�*��aC]����ÄӤu����ULMMzlY�Qq�фn�����`�ɳ�2+}�s������--��q�=8FG���D�m,�E�.,6��ܖ���2�)���'�9�k캡��o]�܇Ji�	j��s�*��D��{���ߟ_<�{θy;�gǲd�.d�R�\��nƍO�>7GuA�y��V��b���4������������i��)A�f�����bוui0�D3�)�:O���V�c������˯v���S^���R��	�޽;
�W����xuy�nC�D��|+{=�p�X���9GG�Y
��жbٔ�/?I�Goۘe�h������x�H]~�})e �J�Fl�W]�_�WG�Z�|/�[�4i��N\�(�Dǫ7�(����!`���a���ȕ��C&�35��r�H�Xb�:��!�V.�>�f��h�O��F�|b�Oj(�mZ�2�J,���'��K}�Q	D�	����-��Ve�������أ��٨檱H���e�<��˵���Q��������G�
 �\z���v&�v0M+W�L�۠�t�5��=~v/9����x�ƍ3+s��Nx�ʜ1�6c�2���׻�Y-`�P=6%`W�3 ���w_���a�u��zwj7���������I)�>zZ]F���硍c�~t�W�.6a1���ዓY ׃7Z~8�}9�ĵ�8O��j<�TE9�g��X��t]���MIV����}Kŋ?���S��l�]�+��/˫tؙ�׃,O(�ȸ��;�4�|@����6¥�WI�VV��9B���H�[<
����m�E�������[�����<��l٪έX�2��M�'n|��8Z�2�;0he�ڝ�)�g��PI�(e0X�b	|�XXy��ץ'��
��3ÂZ�d������)�P� ��>�-=�^�\L�]�/\yk�}kk����'��b_afSU���Uc��w���Y��Y���SK��Rd�����L�h�s׃�� ��3�,�U].�]-Ԧ�!���8�Y�%l�Ĺ����e(��6���1��l�B�dB�I�CE��`�W��b��N<����p��Tk2�,��{=6�$o�g��������}�C����y�����APra���w��YM�U����[��U�},Rr���9�@��ZldL�2Bz͵�����Nא�}6Yq����e�/� -\wJn/�������h��ĕ$)��|Refb��ా<�lW�9�T����`��b'x��}elLu^DvH�4��HՓ�����B]Y�����ò�~��?�z����O�o�d�'�d��(�R"q��AxG�d�#e����U.��i�r�j�_D����,!Sh�6cB�����Ǯ��+4ؓ"���kVsIY 0��}�g��=T�6�7�&��ey�@c��t�*2�����d�0����P�>�ȶ�)�Wa����S{S�,��_��a�?X�Ļ�����O�M�k㊑�\�yf3A�I���仱:$d���W2km�4�U?����c
7I�,����
���F�X~M�,�=��{M�ϯ.��_�W�b.<٘	�&n���j�X@O�88^�K�J����o��'���av��\A.��s1�6��'�s��Qe�jO��K23ղ�+Io5���Hhoui��W�%���j��m)Q��+�~��]3��F�-�����vo���E��mo��T^�0����R_s�U�.�̘���.j{4���9�J�$�O��U=j��|���=����&&��Ls�qzo]������ole�Z�ck��/g�����8�g�H՘�W��E�X���G9\*$���Mb�o;���g5!?����x@�(�Ñ	����L<���4���p���ㄡ���j������g�p���t������#=��g������e?w#��Ka�y�5'���WN��4w��32PL;�֫n���|ã���KҴz�0e�E�IH��ڠqa�^�P�$K�}-���^;q Qm�ʧ4�G&����p�ƽ{�~�	�����Ync��Zs2��c���LoK=M�M�<��k��ﱚ�L���tL�s�S=���Ǖ0��G�����C���0���u��j�዆~��.J
�Z��ү~��QƧ��,�w>�P�+�]��H~cm�u�W���݂�S��zK����*a�ONu�����ui������'�e6^N+���z��d#~���1��^�}nf`v�~݉�{��i�ML�Q�L��ӗ]��Jr��}pP�Dֶ�׭.E1BP̾�:�Cvə���`��w�j�t���n~�����%��i��dTOx��:�V�k���XE�3f�W�U�Xm�I�uNZ�޽�C���V�	��6R�F�ʂ�V�0?� �+ԠQ5e!#�sڠ܀�3�4un����S��@�a��-�w��Q4Bu6��˧!\wD�{�T'̾)F��~�P�ǖ�j��)��)��dg�5�
�+��<SP�g���尟J���%^Z�c������5_'bo,��@#CW��|��'1ʌ������@H5��p��4rxF�^$H��T^S���D��ҥ��W&�M�a���[\��]55%.w�ܗ��,?�أ�؞�u�v��v�wi`�'��1��&)*0i�ʳ�t���	������x������ܧ��-lm�D���^�<t'�S�0��q�J��l"�С��!٧�@�B��i��^um���|^԰t&���n:�߿���Ʋ���q���܌ׇWן��a��b��Ģ����>NY�_i����J8BG�����O�r�ј�/�i,�jxX�쵅�޾L`��PXn���K,^_�|~��xD�-[c���Ox�)����+�>�Ś�^���]�"^���}��5�� �Y߾�U����� V�jh==~�[�DCNK;-�H�&�C�?W�g�:�Ww�+�~]�%k�XEKll�����LK��]ŉ�a��Yd��_��O�JH���:%��'p��մ�@r%�v}¥��P)"U�&�|�/��Q���ø�:�������ZQe�����ӑf����訇�랏��n!�[����Լ���GZ��?̦����' ��
�Y��νZ�s+7k	 ��K(���b��&d���V3�N_<�Y2c�4cKe�kv�b9ܟn�y����sÍ�Do��ʖ¬
]���Ҭ#��XR�n�������iu��'k��k��������]��P*~�s��<��T�9a�i����w���T2lZY�}��Gqs�,4sL��P���#�<7�KO�� \\��Kcm�������D���j�:��^?�5T���~*�1N��Mş|]�\����m�B�">[׏~+tP�~10�����ݫ�p|x��G�y��N9�i��ӵ.88=L�X}Z���\e�M욵�Ϋ�) ��$$�����{ս�H�%ֿ<����ңA�V:*��|)y��$��c������y�.��ERT�{|�(�����j�~����L�܏?�7�c����*k�|�~|����E֬,|�uFr]Ϸ\�マ���WO ��9s#f�lb�?H�����n��9���A�p��E�����ʩ����@<�'�o�W�M�RT�F&^z��N�T��~��O�K!x�~L�M]��x঳φ���~��w_�j������
9K�k���0'�3*�Q��`��p9It�@Q$7\`G�h�1mM$�r5q�'s˜�A�zp�9�M�b�]i�r]��R�Q��;���}�aF�UK=Kӷ��LgaQW�C)�򓳔A��`J�|=Z7�!��d=`��Um!(��v�<[%+��t�f�w�Na����WeE�E}'�Y�W}ks�&�J6=T?���+�U%�[b��EC_|�'\���r��< ��T\�j�!�\�"QOEjrl�bߣ�RT������I ��QG�ˎ� �H�.�u>��/����1�Y:�x<����3��\v��r��4��"/̷�@�Kʟ��璴}�[ꪌ'��.^�ny�>6λ��}���SQ���:��TG�.��I���=������d��K��7�J&���ȕ�c�����N�+���BϾ��a�T�GZo��n��
��e�܇�����>XP1�Th�WB�+S3�
-=F��F���<�}Ƌ<�8d��$�;�� \�}��Tԃ��3�L�WX�F�߹۸��j&tvv�|��^�Ƶ2��t�@r����g�V6����,X[oMvhՈ��W���{V��H�N�>��M��n�vT�2�H��z�A�x�AhO���?�&�-�ŧv0˃k��s oB�ƭ�Y[�gk�%w������f�12��	-:	�1	o���ݡ��Tb���� ����b<������a2�� rk`q���Z ����a�T�éOQ�)��x񚝍M�I�h�F���<�q�fϧ6n	I{��%�ߊ������ɂ#��^3W?��=Aw4û��FC'��5�ܤ(S�����m�2Dz��u�?�)�e�zx|`���g�#���$i}%/�
�WI]r��t̾M��	��N!�s/����񉉹��&b����>cs��4O�63L���gq�3��~�<;$
wF��6o@���{]���'r�����}CR���/��Y

sR9��KV�d�z����"�p�P�HDK��'Y��H�ƭ�b4������s����[J�)�9M�D�?y�c���,��7�t|�:v��O$�����b|���n�gu`��Q	��b��4Z9�f!�@s�Ҋh�X��Z�q/c���xo,��K]L����*��~�w�����T@�.Ү�-�du%#֣�q�F�o�6����H����-����sL8B5!�$��93�9u!K%ޅ��!����ϯ����?�ʱ����[��'��#Ezm�;7���vp}�Ϡc�y�'f�9V���p�ḫ�7�*=�lNm(mi�Q����6Oi�z��O.�m�iT�*[ed��1�Y��w�p��}2�ߒz�Ӊ��P�a��}�Hz���@�8`kkR�}���/B����M�'#+JΒ	%LAe!^����샴ӑ@�Ŧ���W�9�?��b�J�p��_�R�����p݆�ۨ��̓�(~�Z���B7�>ĥ�0���]:��n�{����ٱ���I��E�?��>z���lg��L9r$��͊�d��Vq�&�f�K��*Aa.�2�2��
���[r�������>����٨�E��)����0�ơ�ڧ�auڵ�9+z��C{QT^a\<<rY��D;�y;60$�X�*���!b�F���M�P-W��U�����>��o��%$�~��[̘vK�ya�=A��?<I�=�5��E�j���Ɯ�G�Y����w0�����䢋������x�����f�БdIS�3A+@��Rڴ^�<�`N�k�8t��v"o�WK��aA�c�,��Τ��~E�����z��j��! ����������1�|4�SD5]�v���m!�n���{��*�P������?J�0�]FFF���{�������S0��G��o�_��贲�r@Wz@�;�c�<a�G��
/XP�66Ff�Ú~�-��5��vsJ�L�X��;���T|G�UĮ/mm|�
�:؜x��G9��g2��y�~8���ҫ�E<5��
|ܕ�)M�'�6I[0"��N�E�T7h����oq��u�~H��;�}�X��gx�$���j�h5%.,�8#P-/BB������J����[�,⑀��;Ԑ�3d�<��c�Ζ�}E*EvQK|��*¬=�Zj�k�=�Yj5�����[��U�/I�%���M3���wI��q�ԅ5��=}�~~@bF&+�'�l#$e*�^�]dɞ�G���H� �;�$�@�x�
����ٚ�S�2ngc�wY��Y	���q�9M�uV\k�]���l�t�h�1�-b��I� ��O�e�ӟa�nO�z�Ɠ_�M���Sҕ�!�r�#��4����q�%����%��j��T�ii�M��	��'�%$�U�N�L�O�|5椫����E��ˋ$;�.�D|������M���ˏ����1Qݳid�Ш[�{�d�u:�Q%
��\�*dfM���1�z��ߕM?�"8~�!�����>�9���80�����lUy�ؘc���oi�Qڧ����B Aj޺�� �<_�a���?�^L�Tl�\���Y����(�K��)I$Kï��_[)	X���`�ّ߿�*���m��}��C���w�b=��૮�1Jp����*��Cg+� �T�P�l��>.ƃ��%�.����]���7I��a�����ؿ��37}7�;���
H�|�����z�}S���2��8���W��c��洹44B,U��_�^����� P����b����[�	'�z� c��x
��H,�V��R���5���+��wQ� 9�U����}`�P9���Z�i�p�	g&�8^��)h�'B#�ԋ�Z�+�x�� D���*T֗!�H�%A�ǥMO'D�Ơ8���z�q}�M�3>tR��d���vV�V��j�(d}�e�d�Z��=�|�f|ֆ�A���{~�}�����@l�C��R�G�s�i�0j�_U��H��d�x����
v5N�..�9  ]A�mC>����l ����ۤ�Z�ѕ��ڡ�|5�x�x�s/}*��7CaiL�x̛_H;`�u���Z��3����P�h�������/�<�5v�v�����dL ]��
h���+Ԯ�1��fE���� fm����]evw�}4�zoү��*a"TO�x�xW��l�7MS0.��f�ڀ�z��c¢�̱�g�Z%��*��ޠ+I�DbbːrDzs�r�&�P���!�����5\�v2���q�p-���	!'CQl\��q����IUWi������v��3[G���fe��9u�MD�e�g����g���80�_���tP�MOO�O���]�;N�&��XS}f����\��f��4�v�J��rr�P\J)w��nDw��+��G��&<���zW�<d)�|��)��+髧ix��f�S?W����� ��j�����jp���h5�"o/{�Je/��4��;���>X!p`��h7�®c���D+�>��U��5 [��=���7C��h<����E[SS����=n����h��Y�v�;B����ǿW3�[��6&mװ"��#�۾R�Cx��zo�8���!�lY?}��^�^hr^^�����R����
?U�Μd�h5�/q�/��n�r �F�2q"�1�?��cW@ +7˽C�ob�mgdH��w�P��6/��#�D�|�ؕۤ?�\�M��h��ߍ���R(��s2L}��^}��-�q��Q.�g�bR�Sy���� ���~:��^r4�ۍ��+5~Ǐi�թ�VN����/~��j��	���/���4g����"|�,����ڴ8���n�guq�?6�����Pl���"��+Q�I�~�^��A�E�6ϕ�5��o7�z��e��l�ף:��S}�:R5%�!���u-�z����N1!0�h`r8����?5^Q�����ԣ\������J�z��xC�0� E��߿3��%C�@vӺu8�����T�˾��k�BnվT!�0n)?��9��K���zHX_��a;����*��۽{�U��"�{����Y���^~�bS�
r/Y��Պ�:���*�?B����N��b����t�Wy�
R<��}��� ���5tt���Y;�I��tl�T�/˭R�|�˱�:X�IQ}�t��d�ӧ�z�4����&)c��J����[K��b�Ch�����~��H_�)�\vc�D.�BIs��XP�K�Y���3ͥ6z�u�H���|uuY	����9|��h���
r33�Z��%��v�*]<0o@L�͚nmC����j�4���F���*�I���f	��ق?����8��{�ȏ����Cn��{C��Y�Ə9�v�y;E<F�O` �6�ƍH&�÷��w��AnW�e�nP�|ޟbZ����b
QNg���Jئvn���_JѨv(��*�(�. ��5��ojL��pa>��~1�q��ߋ�����G$tAB�J�h�Gp�F��&�~�<�7}w|/��Z�f&�e� ��2�)20V��iOs�o��wpJ�*�;�����R=�(���&�ݓ,���t~w"��*[��%�vZQQ��h[(oe0J��dTV��������G����u[�fꗪ���w�O:����0a���v,���KC4
s�@� C�)��Q�N'Vo�V&5�G���w���|�������\;Z�@u��k��Mcu͟P[����S������pᇿm_�}�!���iȣ�kZ��w�E���Mc���J���q�}�f�
��������Jf��ع�8��^��A�����9iq{+�4��F����l�K��� Uޯ]79��Ḣ�3�Y|(+ �w��6�f��u''~���t�/�ݲ����_ׂ��Pr~��~d�V4�B��l ]���ֆ��D5n|*˖��9�}���j��p#��饉�������'�L(g���.�0��~::�,@�Wep�?W%��D@�7VB�?@��S*��7n	�ӎ*ۓ�5Ҝ�t�X��������2�H��2B_�Y��)�SC�ɱ��?����eڻW��iP`ŗX�,�I\OѸ5��}�֯��P��e˻n���$�H�ʳ"�#~J�t�1�> ,9��F�t�����(�s!�Wh�U�[�F+�~9((:�#:..��Ai+���8�^ �js��_.)
�P�Ɖ9��ޛ�Zb���v1��K��>�]#{��0� �/w�RMAnɺ���%j[|�y��N�����Z}�m(�����m@AȌ��?�h.���u k�����A��S���n�{��#蝻5�=�1���[��E�T���qT��!��v�g6�� ?�y�'���ύ�o��ǝ�n5�P׉T$��X��y�L��v>nyy����;�TMA��������`���Ӧ1���No=�3�"�˺�W�@.��G߿}�w��//o�q���ڙHUL[	6>�܁�>b ���Wm�D�a3$X͍#s E���K7�Y�����Ի���U���^_�8�y��]^O�Wk��NA[XX����}�`R3
��=�N�:�[��&�����ML�����ѝ	����b/�g���>4[ �};2�(�,���?b�+�P���
��Ǿ�xG@$�C�v|�&11LЬ{��3sGU�?�A8�9(I궃|�_�亜����/o��HzpwjH��Έ�I�g�-��>8�P�d��D��[b{���~_"��C��@�:'k�����`rٖ;��G����B��K�Ɉ2��w�옝��1�;<	�N�H���y+TԶ�u۟8x����95T�g��1 O�'��T��ظV�䏺+O�>�&�>���Y�s��~��w����G�>~�� �3;ʹ�y��X�_a4���&�
�\�1�shn�|��I���
F�AT��Rxa1�������y��P]�%�����/�\��rJrH�H���=�����ii�<\i�A�-xGP�&��"��훦���)d�ó=���n�!�����!��[�֍�.-5�p��[��U��d�F�wF݇��UTUl;�B�BPh4�6��C��׆뀫|��ԙ7��w�&���a�6��&�$')c1 �"�m}TQ�#��PO8ؓ������ u������u<�~]A,�w7�q(V�	�G&�_���C��%��A�'�*bJu��6�B~BX欼����]ʬ���]�D������[���&��jz�N���;�6R��Z��*e�n���/��ǵ�|W��*��Y뵴ҥn����.[�Wb;|7��T���t^�ء:���5��r�~nt�-uP�I�ۯ�菞x�M.Q_�s���t5N��E�V�h�{@�%�V�n��$u[^K[����Mo�%C�B�F��t%�3/.h����J��R�8����|�8�����J����3CR�a�ҝ�Y0��_�D���t[(k�J�����L�Ȼ(�l���w�U��<k [�S��]�4ӛ��b��,��t���/8i����S?��ڳi��&+�c��|`3�|�ji���.��v��<����j��	����ͣXMC��7��6�X(�B�wf9j�R10a��!�缵]��&��!yZ��j�zl>t2�s�X��H:��O!8�6:�%���P% S�^�L�?qq�\���v_v�df��F�pI�`ie/��ΘA�n��Sa�%f��5�zz��}.���W��|?J#f����9�|����(1Ӄ��V�Q��y���+��V�C:�ĭqî\�pj��p���2�t@2�8���$q.��8^]^�hX�ѧ��W�F�����]�-�θ�k����z����Y��4�~C����)��ު�-\�G�F��r�AȦW@���[�G̈́����X�8Χѷ%�4��d��m�p	���=!���^�^�,�oE(X��_V7	���2-9v*�����{�o'�㨾�¹�[Ӽ�a�e;��?�}������
<���:��>��ޯ�:,�8�D� ��b��u»;�b��W,�;u?״Y^�wB.Nnu�Q���l^�ZA�33mҹ���C�k��ZA���֝��xȷ�{�߃�����_���!q�Ǯһ�'ۘt5���S���]�� �4|	�j�*� �>õ����8?h����Be�b��Vp��eg��Y��_��3�R929T*�:��	�c)db�$C�T��:\����R�g�r�m�/ɋ�0�,	S���g�K����aÊ2�������*?)֪B���;C�$w��@x	��x��%�R̋W�J��P��H�v�{]����>�?v���͵%R~�56K�������o��W�K矐�Wg� e�t��m��Ʌz��������]:����x*�;L~�LiU�Q���C���6�c�L�o����6���� ���#>_8��}�Y��ȡ��ag���T~%,U��Qz�E��`�xT?��,�-�v��Y�x�MZ��5��T�	�M��+@��y�]6���Ҿ��[1�6���ݽX���x�:,G�.��x ��P�Sn�9����Yt�>�`�yăW���|XO���.�����o��g�b�1��,wm��y�|�C_�Xj,�ʋ'K�۴-����l��񭝫xJ����t��v"�g;��G���DE����Z�0K����"���� A�=��_�zWT���o�u`�jC~?��_��=����{�߃���� �MK��i"w�ʝ����ɷԺS���N���8�0mzs˥י�q(�n䙂Τ�8D�Z�6ð�"�Nn�����'�rv�y��-5n��XQ6Oʸ�x�WM��<Z����
�[ا�໾\�x���(d�3{=��k�k(�s��&�2�Ѥ��Q�!Lk����o����`(���C��KW��ޏ>.�Z��X���W(��~3��;�]f��ϲ�?�`���	ʚ���>������`�Z=xD�4YN�+UK���{S��=ie(���n֕}O��3�幑��5��|�:�2�����F�J=��g���a�(��~fU�I$ ��]��r|�e�t�()�o�d��e�|m���ú��s�m�rNi�����fR���WH��b�����Bf��(�Y��C�[�z�N�}~�%�.Rj��G��6A�RY�Ae�N��¥� .�S�M�什~�?pa��&�7�I�̥;ϻ�l��d���]��/vc�K'�3W��~7	CJO^8�[�ላ(%U�z-7�Z�Q���9^Ct�����Y�:�Js%���܌O�\��v�s����Åǩ�/V���Syq���d<�yN��[�_OfЪ�*s���vU������(�µ[��S��~E�!~�ɒt�����:^�2A�gbL\W�VZw}�������3������]
��7&`sO�Q"E��o	��Fh�yO�m��k ��D�J�����<�+��rK�����+���$3�M�Q��w۶l�K6 c�H,��+9gk�Q1��v�(�M4d�᯷�p�>'���P��Z�i;��&;7�.W�wc��b�C�$3C���|��	�v�(Cw��h������i�Z=�ɝ(��L�l4��T��h�]�+p�$W<z<�*$�:2�/P^~&/��
n�/Z�0<\��/��?˼1ͬ������ J�T)ɀMX���bʩaB�@�����H���hY�E�J	�
�EW�x�FJV��m�~8��h�=�1�J=*=u��R��p��\.N���._��[���IPS9G�{��O��h��q}�0P����V;U������{�5���� 8��6�� EA��X(J��� ҋt$��Rt����P�I*����W�% - ��I��s������ˋd��S�羟��vg����+Y�����F=��!^t�ߖ3��A��S3~�FFد65~,r�)�O��O	1Đ��q%+�U~���G��ǻ&i)��²,�+rX\�{���oTX�\~U~g�M�3�lM���r�At�{�7{��wDȄA���G��GђS~�S���]���mq;�]H9�A�8v	f9^I�1�WO^RZ�<�bs��\���\��?e���� ��:b�S�YB���wO�k�◉=�)0���n�K�Q��S��̉�J"��YI��C-S��6�Q��D��z'���Y�������,6*EN@m�g"����N�os�N1�]w��yY��օ��ܯ{1�a`YR��d!�]�R����	�~�V�ｇd-���_uLl��+1��A�x?P���E7�kװe������g����w�k]�A^���)˻a]�����h�fo�Ж}���&����h���W��-eT�rN��0+ߟ9^#��1r���vCo�B�]���T���&����:�f���K��ߨ�����K�~2G��>�"w\�~��㕡���ܨ���G�$�t�7?��g#%r/��+-G1j�=��f1��B7��E���#�Eϴv�&_ύ���XHm;�/T�čs_s>�1 MkTt�l�-��y�lta�\��\ ��q28�1Ja^��V���l��c-��1AoB��9�9��{���I ��.��q/�ιj3��Fol�|�)�y.B���P�է��.!p��xSc�ZĘ�¯�g0k�J�����n����[�Sw��<�Tk��f�W��y;"l#'���h �W���$�J��nƐb�S;��H��DSBɯ�_��C!J+˞�W��:�E����	���*r:���<k�༦&�w�y���Ǯ+�!�O�%�m��U��k4)�D�.�1
�b��3��ϵ�'}Zλ��I��c�&?�t%M���bD�3�2�}%{2��ʰjsi��y��S��eՊ�Q-�<����Q���a�X����>�O�]���..V��� �������m�A�9߅��,f�}Km\%ѵL��'�"���z1bw��ظ�둟n�uO��d�!	�7�[���۴3��������핪�ɫ�T�=�ZQ�G�kU�a�غ�ۃ�לB�J�l������:�M�JsH������<!��5$ka�<vc}�k}iBU��U���:��Q: �O��);%�k���a^ZŲ�'ri���}g��=M:�d|���~��	�G��q%���!�N�m���e�4ks}�LVRS��jֵ�F�x%zfﰖw�p��}�Ő8�!x�8z9�C���)��H���<,�N5_���}�U���Z�{f�1_��Y=��Kм�(�Ŝ�؏���"!��~_��9�`ۃ�;���z>�K�J�v���~�UFEԅ�Y+v��Z�e�X�;����4��$�/�ߝ��1���`{���E���Ыv��~���&Ԍ�4*m�?�pBz)����
M�*$�!���0����/-H�tۛߋ3j����ƞ�Zۦ�5���ݧa������?x߆��ٿ7"Y#�t�WZ �TFX��������;\f��mB�i��ά�}eg�}1�?�L�>��P{x��n7��M�#K:5f�qB��m����xr"� &8{g�L��i�e���{�u@0宁���jGƐD���֧'T��'ϴ�J�?�=�{9LJ�jԀ�a�T�> ��g�C�L�WN�;^ñ0��J���L��ĸU&�W�K�Q�ta�
)�Z�s�C��3[�G{�9�9#R�6lZ���~��s��ٵ��c��{�T���W9C8����ɛ��z���bo�(I$c h�,��YmS .�90�d����9>g��j�k�3�N�^�N������ʩ;���٣&m�F��t�G���j�6���'���n�U�G���q���'rșLǶ��"��O���;la�j�b��F4��An��Թ��p8�poq���e`����}�Op��*q#�?�6���wP6ZOJN�Yj`��L�V��H��6�����˞8v|y٬�>'��p��ed�i����f�P��Y0�:��¸⎠�3�����ϗ=����J:�
��a��w���eh�������aʲv)e�3Y�Nt�]y'�ʩK�\�rىB�tC=�4r:O_hUY�)�xJ(pE&Pj��8�U�z'b0��V �C����p��%��~@��l�Q�]1�o|u�1�?��j{>(�@�D����e������|��ayT����/z���U����zc�L�L����F]<�;X���xt��a������"3]y"|*-��%Cr����'p0�H��MkiP��%А���"���y���\ۊ���U�/�.��|=���5��J�CS��j���q�]�q�k>m��%i�<L~^�ȼ����/��L��w�'z4��r21@�lMV�w����#s�}����:R3�D���*�ڵ��ڱm��N�1�on��~��.Rv7��)�;�[<���r��D�	�+s%ش�_�&r2"��H j��d��\���^"y���Q�8�b���F�ԟ��[�y���˾=\8R(��AvM!MU
���K#�5��K���9YiE함�tf�}�K��,�F�@���O�Y
�R���T	�4�Ijs�	�u~�)<i[k�^\���P�������n�2���a���.
Q��V�Z�Yk^gč�M����C���N���p[]y7���}N�_���������b[-��\qK}��2Q����s�]���<����yW�[�es ��i7�GM��i��@�'��(O_�CN�n���K��T�Y<�����}��]Ŷ�<�=�&�R�"w�4�,�c��wN>9���40+��S��WY�m���٧V�5?�ޢ�0��.��₞+Gc��Y���V���*s[ɥӬ����X�&�^�1�J ,<}@�Y����П��&>�u^�5�G�zo�<�]8ϩV^�4���`^�aEP7������mR�����M��������[OM74�V�eq�q�w��3PI�[���l�~k�m��p��+v��͸�ɹS����������ͬ�A���@��n/?��=O��ݣ��A����K�����Xk�F��/�I�=V9���.���p/��y���7.�)Ё��u8�3��Jf`��������_����C$��1T�3/����0�\C� j��u�}���p�	>�w(�"}��&'f-��H�`�*�\�_�|�?񽁒�W�y�d��*&6��?�!��#�d��f��έ�h�Տ��\�����=�ִ��1��Y�X��C&F�U��&�>�/���x�	\z�o���U֑��u�'���O2��^�yo*�W�FP{<mz�n��͘2&Þ������������}�{y�?�{�n?�u����2���x�zU̿oV/��(�#W@������Z.���k�xPp���&ɸ�ԡ��`b`�~��Z\�f��G�9_�����ư³�R&�*��iκE�6��JY�D�\J/�-���o�)W�Ǉ�~㱳F(_�?S�8.qi�a���É/�K�=�6�x0����m=��}�|�T���(&<��N$8�/�"��{�!�7�BI�
��_m�h�N�s�0����J��ª��*$x#I��2��~�T��s������n������2�g�,�œ�I�C�b�TVK	�b���fL��A��/�s�Od"}A��A.W�9�)=l���_9@��P�8���^s��C~�sF)��ԽC���ϧKg��5��<=yɰ�����9E����[�%Uo�︜���Nt�?�v�<'�m����+J��웤!�|{ƌ+z=�\R�`�=�mʫy���}]�rȑ�����F� ����ض&��q��GXg�y���
���N�0p����t��9�X��E������'�9tx<P�}1*�7���S���]uٹ��4H�p�����]�N�Jr��Gm�D��&�J�bn|�@�c�ɾ=������Ơ3f���%�!f�E�%�i����xM ��z7�f�k������R-�
{��XP�*��dnO8Y�$B���}��?E0����f�"N���&�?���XX}�[3L���v.�k`�lND^�nL�B�V��-�:������u-Ruو�f �J,1ї�ced`�������{6�,ّ�%��P>�P�G���;�b׾���&�@#Ha���(�.L�xzۛg|"�fn3G��=���h��| ��V����%3E˹�I�$'a23��;�w���󂣖ɥri,��}�T�ln���J�[�BY׵�=�+�ϷD���y�в�5��G]Gy��X�ȱ�����w���E�vW����Զ�
??�����}@P��=��C�e���]&Et ���]��an�ݓ�Aq��:c.r"C���b��P��w�d��٢���.g�]�RV�+�
�{�黍g��6�8��7�j�D��-N�c�+��9��>q�2�:�ߝ�7A��Y�|7��s�^����˵�l�����IY�@�.� {��Kr�������`�{�+F��M�{�>��'}�+�Pàn`�f`�h�
(����77=��$���'\���*�D�����M�ۡ�u��G�H��(͌���r���LL�rHa��o�w�l�;ڦ����mj��v��^�k�	=��=&�b�IS��S��h��~�ș��J�?���mH�Wu�U��~���gp3h/�����a?6�Fk牳����{Z鈳i0 �����H�9����-�n�u���7��`���R4�ٍvQ4ٻԲ�Nw<!T�_o�P9Հk;���l0���۵<>�71�R��P�� [��BD���ͳ[-�u��7�)���Ώ6	�	�S�2�W��2��o~Uk�ho=V��?Fd�0ݥ�;_���� l�Wa�vzX!��\�����"�A��n�̤�:�-�s`��/'��'��\N��'pJX(����w�t�;�'X���M�,���*.�1=iUn~n�Z��?)X}a�|s+��i|}�1[,Ho	�
����-������"QR��Ak�W��a�s�{1�e+�)�p�g�mC�[C}Axt��$8K��V2p�Y�������a6���0��}�9�V��t)?#rl��ն�V����Qe�T� ��G� �_9͘�M��g�Wٶ$ήR��Е�LJ�Z&�l��	\���SW%���= p���~8߆�aaPس��4N̴��g�@���h$ȡ'w��8Ə.<;jwT�BK��|a[��H	׌dK��J|�c�ů�Ծ��+i��u����I��Z�e`H \_x�4|�k^���.>b�S��-����|��W�Ƒ��0���LÝ,�J��5C���u�\n��s�T����=��h4��Z�Y���Ч��}<쳪�ֶ7W0#����?�ڟz�b&�,���&�ڗ/_�
��<P:5�%��i�O��?�(��lK��ox
�/��t)S��@�U4mj���ާ�P`�8�Z����g���ÿ������+�^�Y�\ؘ7��Qf��"c��=���O����v���]a����N�~]���n�l^�Bk��Pdd
�#���qU�99��M�#.��̯�|�z��+�}���R���D��&^�Ŗ�9LU���L��X��5u��|� �����H�AW��"�ԩS�)Ĺ9�USl����_�i�P�iFGG'U� (k����gt�RR�J�EQ�mmmZ�V�\`�Z�lyg`�l����7��yF~��d������ΘĮ�������b]jj`����v�l�_o��]YU�gddt��_/>t\�����']`��Q���M�=�L��oD4_���p'W�} �W����m1^E�B?�����_�F6��c/�2�/KKg�U�<�[\��6��Hn�@��s�\r~})�w)ʯ�L�]���������ݵ��x�l��
�ui��)��K�o��T��^xD�M%���r��602/u���*@�� �[ifv>>>Q���L6}�c���}�h�N��R4>榩8sKG~5�9\ Bq�,�2���шZޚ+�!��f�5p��G�W��^��Z��e����]�=Z���oB�=����Q�S,�F�7-����G�.p����Iex�I�;,���@{"�NM�	�Ƈ�L�f������d�$vga�XwZ���i5����gCCC�ee�sz-��1f$&%��/�9�h:���(9ݏ���!ʤۮ �0��kdA���������T��,&RN���lf�+%��Б�2�����mu�[+P���b�_�>�e�f�{m�c�pb�J���Jt���[��/A��T�­+�=v�T2��o�`�\Y7�� �v��@�Sݏ�����,�[s��9}�a܎��>%��q��C-�kR���yӶ��X��J�Dm �<�	�e�����[Ri�ߣ�KyF5y~����E"�g�R%y�'�o�A��Y`���� �0���۲���������<+�Sݪ�uK��I(�KKA���l���*��ќ�2�� H��C��!'. �z}�S)����h�v6�5kWf�۳�g��� 5�
zB��7�O.҈�k��<��T�^�s����O]5#h��|���>4]'
�4	�iA���9 p���h�����q�'\��Û,����}��X�,ɡ:�,/��F��Gi��Zp��]Se"���Y�)]�ņ5���>w{��p��w$�D��ޜhn���G���`�f�f?%_���۰]1�����?�r˩?Vɛ���lW�;/��5X�A:�r�L��˨��Jk��|��ڍo�5�%�s̖2�R�n���'cM]��*�B��[�H�wzJ���͔@9,�>Q��ͨf�3�z�a��u��w%�I~W���Sc�6��~8h����� ��`�*/��t����=f ���c��M�~�}������x�����һQ�n<����[O�L�n�	�ǒ�?���vU�4g�b��K�)�\2��ތR�$3w����=>�D=��J�D���iM�-�iv7C�%�fU�e���v��?�.���-��������҅.�hw�s�:c@uE�E��RGGF<k^W�Ǹ�`�� //�B�5�!���۪��H���P��pS��gо���Q(�83�[E$/)+F'_ߍ��7n�஌�*����w~��� ��p���)B���j��R�+��k�.% L�<�Q),eN]�uD��-�kR�Vc8`h2�?r�.��&�0�9��D!EQ����t���5��"ŏ�Y����%�������M���;��	H؜�'l�P������l%n�	g�:$�=�Sd �kg���B�Tm<r*M D�y,�Y#����>ϥ���%�0��
�ݥg�Y�������sa2j�J��U.�@�ֹ�cz�s�S������m<z�T�ұ�3��u������-�E��h�Oc
�j��X?�1�|�.�� ��$v��ڙw��(	vHT/}��,6��Ʉ"}��-ݚ�ҪP�W���lF(�x\ڋ o�{��k�$��-��5uxX�{T��o}��L)�]A��Y���;G�G��(�Ӈ�w�?4�����͆w�^:m1j��������K-�Εԍjo��F�f���t@���F��?gW7^�E�s��D8(�=:U��[I�}���G"��#@�ν+n�CP���μ�z~�jW����ڭ��=S�s������gE]�6��q�����T�������쮈�Zl�qqI_��;�)�J�Վ�������2C� ����݉�����	�{���M*)�*y�M�[?�)��[��E@-�7wŨ��5�:�]���%�QC�V����ms��� e
e���Q�;~|c��O�y�9o:b�A7�'9�A@�6a��S *�ox4�<�'��mʾT;v����5܉��7��פ����ռ3695�5>>.���J"�o�n��qRq#{��V�q��*u�N��Z�XDH׬�u���+	x3�ت|�L~�`������/'U�EsH%�VW�����@/��I�J;8��~�Ў0x�-b| ��:Ǯ���	@�*ǔ��H�$n�j��{Fyi�3KjQY)��ȏ?n.s�D�Me��������ڝ-�i��%Ƚ�������Q�8
�IB�72x�+ng}5��:3���cW�-V�W����ȋ�yȴ/6%� �ِ?9�<��ߨhۻ�hX����6�|Z�R�2nW������0��i%D����O��L&��s���������.�Cp���WZ�О�2��h�ll�n|+��i��E�'�Y�Y5��\T^�m�zK���*��n�B����;�&���p�G�f�
��ᨆ�S�#�f]�M=�{��O��k��4�,^TTL��ai��*cr�ߕO�X�eɊ[�C*�n6"���l<v�a�v��c����~o�]��Լ
�zp�ޡ��~g,3C�����R=�7��
��k>Ԭ����Oi�h�F׬R��3y��_�n�Ta?�5f #��L	��Y��GCFF�
����	���F��bT�z�^�� 
�BJˡB�*紂�.�F\��UJ]�?�`��[���`��GO�
�\Qjj<��9�}e���f ��G�`�B���\}��l�\TTt<.'_0�jv�{Cv삙��a�Fnt����Z�;�i����U�B��\���VӅ�KQ	Pפb�.�a��gv���l��:���zi&�'��]��4�t��m�܁�\�
��{��;����\��sEQ(g����K��{�(!?��И}V ��0�Z;0s&�j5�������v{��+�@�{�W�䝕@�h���opD/��I�wft: ]7�kdǍ�W��-!�)�.�&�wĔ�G�ݜ� @���jݡ}Sl����ޛJ�S�6xr� 8B]u�P���������i`�ܩ_]9/��:�t(!j��9/Be�/�6g::�������5/�+b.]W�,��T�?pojLRf�Ϻ/${걺�$����=�ӡy�� ?A��e��z��W�ה��8!,d�]�A��,u�2R>yM���#��P���0HL��K�Ml��S���wܱѭ;��ԩ4x���f�-yH�r�3�n����+=m9w�x?@�JGgPP~���n蟥>w�-�+&yQ<��$����s�z�_�PfX�z2�N\�kg�1�WD��Eyq�T��!7Y��`��
��ܣ����
¯i5�<lJ�G|�UH��	�&*�n�(� j��ChK5�_�5]����VWB��Q�ą��/���o�[�A�����%ƩD!;3ڡ���E_�Wb�tn`�]��Ǐ�>�###�8;+�.Ι��������·[� �j��S�=!�U@���_�f������V+��8��j}Q;��T�cP��)י]�S�	+��,�@� 7&; *�
ei���9v�
���j꣔g�;���ęJ�H�R�\Ks�1�ąM`�Dhʽ)+� ��F&�;lƿ�|�o�
%ˎM�ߧ|���t����W��w���3�jˢ�g~F��<;�5����|�� :,^�7�~\���F�5��p�&���.{���f�3�a�-Qqs+
�H�d��5�j��
�>��`c��m�+o_�0	ʨ��ni�K/S�?sE ����:7UͺƳjj����y1)���V�,��Y��٨�RRR{�ϨE�{PAz�?�<��P���D�X�#�(��q��;QMI���v�� �X�ڂv��� -��j��w�-�җ?���K����rF�sY���_i��n�\�ڷ���u7�w?��I��[�~���t��1���݅�v�V;��P�?�_�ԹT����M&�(�E,�"y��w��E��U6�� 4�ȱk�{0k8Q����V#�����WεE�5Z��W3R��ڛ��_�^�
7n:u�/ �R>2"lj|k��쨤h���b� ؜QSb?�v5 ��>��;&����x�~A;ِ	�S�~4�}�C���@�sG;��э�PcGǝ���35�]-����ӻg��я��a�;��{����ƚ7�<� �#��m��fo��tDTTvEE�PHbé�����h�C�e��掑���;���2��ўZX�2�7����ٳ@�NL�q�6��rU5���c]x�~�2�'���l�b��镋ўk9�M<2-5�bMr��e���Jƛ�>������˒���y�J����9O�Y��ȞW`��!��Q����Z��_��;�ʁ4/�S5L����{�1mȷu�8��]�"�S


/���%����>��m?G��5�}o��Js�H�SƮ���:���?��ey��̦�.0~���I\�����ɩ�����78b����hk+����F"��*��cV���HRRa���?���%�� ���t��h���$�:��H�������Z$9wWJ/��\{�G�+j	v�d�� ���*g�غv鞿j��*�h����V�@�8Ea*ٳ�gu��?6�n�O�O�;::�f�e��w7��6b
�Y-��G���C��	��v����x��K�n��UU�vɯoN$����kG��~� A� �Ĕ1;[[�;��;�T��ʤn��'����ʺr�F�X׫:���x���tΟd�������.��~�{l��l�=��$�����ҿ]I�U���&�̉~��V�9���^������`R1uS\�����x����fff�Ǯ���L���"18y��4"��.M������%���ˁ����)f�X_�ߪ���9PZR���<?����[���YS�4
o���;;?���q�M�8�̧׋T�y$;8:�?;̫���P��h�ԥ5�F������|��w{?��������՚)9�\������Lܕ���EFR��/��z�鎂"v�H�����z{{��mm'��2.;ű�D?���TSS�a��ID�FNrh���0��_&�3�)�����9�[T��\~�~e�A�������ճ�6�<�X\�� ��������~��+++*�^�S����k����b���]����[���dx{{g����`�����/_ڧ��E��ʿ211�E���}�c������"��! m��;����&��I�Y\��ot\eP�����\Gg�+��x�G;x06�aø������Zz&_�&V�Ԩ���H�;��S�H������1���%�����]�Ȉ岴����h��c��ס�\���Y��㳓!�Ԩ1�����f�/jd��>��N pE�NqswX�O���.LMoz�|,v$�	m�A��"v ��YI�P薔�f֨��M��I�!�
���Y�m}�"'�$���������ynq���ak�Q�_���p��WLe�����hhh4�s�u�UL�NPH����O�P��ˠ6v���FS� �;������I
�K�`���x���mY�hSɃj7m��7o�\��R<��;���NO�`�LC��
����e _�D��S��h�-��Q�y�NIRA!�}��*RSS���j��aB|��3g�8��9!*?�1�C����F`��Й �9�:9P���|�PҠ���.�2�� z���O���p&�u	�o��k�������������
�-�@�ONN�Y����cgg�+b��5�u�1��\���������;��AR�	�A���ZZZ��`�F0>���5%9�Bw�a0�\�⨧בI��_������`��~� ���x�,�XzJ��";�\jw�P���!z��ӕ�(��"oaA�X�򢉟��'ii4��8=Y��f>{���&sy�%KG{����>د-�~��TQK8�2ޟ�VqE�.�m�&t�(�߳5����_U�$��` �%��Ɋ�8A�5t���S����z��������;0��a��f��pC��a��� ��l5�F�>�3/�� ��,A�D?��S�W� �����H8V��<��� ��CI�U�������YM	mO�'����ǐi������[��qq,�9�۟�Ė��e�(��k�7<����Q�,g���|�+Ն�����{����ERJJ�_d<���秅@S�r�T��1�2�&45��&4A^���i��qE|���#P"/_��*++��b___T�$7�`���6-��� ��(b�Q+�JK�, �c�F��cK���2����;r�K��F��B�_��'6_���� R����I�UU�����EA�ei�ȭ|4����Y�봋���tZr� P�M�<�&�r.l~&�"���)���&&�v�/��Y��3�
���_�x߿�1=�0!M	��������|�xh]�Ǳ�.�x�v�'qtO?mJ�-�|rH����9�RuQ��)�!�+PM=�����1���h�kl��4��uS� ��#�\\���q�c�y:�Yԡv9����B����e��`0��JO�|�Q�����+���k H��O�@�h5܄�+��Ç0�?��NHK���jS9Li��)�Oq��Y���w�q|a���p��R�{sNP�i����� �g|���:�CE�\Md�g��]���0{Q���V��)�s�da���vU���u'� �XF=?5%�����+�侥�A� ��MZ����
:k�=�i���!t���H�R

��5qo<� a|��4 &n�@$J��w�Ґ7莰ބ&����ؒ��� \�;���6�6����X���ل������ƺ���'$$X��j'�=�#k�_���*y0�cZ�ӧO�����D��uv�~q*�Y�-ѡ��$J��sss�-���;�yM�Q2�BM�FFF�>���q��b��u�-���n	xp;(�M榦�� ����~��3!���.>,�ԧNA��b��=��W�X��'< ȫ-����a�!�
�
�"���Է�xyy_��l���䢣���> � @귾�Zd_��/x�˩�j����vJJqN����mG���~b�X}��R{o��ϸHuk㧮���r��B&�i�����(�4:#���=ҺR������~'����3l��b1H l`�b��c�^��s�:Н¾���ﻎ��TF��^��Q����m͚r@�@����<��h�eē����.����*�~�aB@A��EM�4����p��*9ɀ���D�Sp�83�A�r�Y:v�lo\�s.�ڲ��7.���Z�V��IP�='�6!*�ӕ���M��*s@8�W%@��Y������\d)�5d=��jVu���ŋK+�����\�j�(B��^__�z�uĊ��|��['}B�����w:`���
��Q �\��L a_�-�*��]bR�ޤ�� ݀Y���QO04^�V�z����XZ�������K������P��O#�?��%4%�~�ɼ� \㯱NɣBw
��~��v����X���m����F��m���;�Φq����� ��K�ݤ���oV
.�z�-%�߯^�� �.J�ռ߮OVi�n5��j\��J�,���&�ӪDB���}�	�d�U;!~�3�x�E�#q�kk���� {�}��fT� Tt�N����g�DMZ�ݞW��ߋ��M�6�]��
�P���њ�[��6`��K�ѿEoU�QŔ�]�c(�b�iaT������{[EM��iS���^�����U0�ʗ�Z �`;�N?�����^��ɓ�j=�su� lTy�ed��靉p��ē���e���L�Nk�DW�ŷ�j&�Љ�3�)Obo���N%{�F|������I$��N�WC����-ܐ��)��^0�o���MP]�6�s�hR��4��-j �`��4���;FO�N�n�3����(�3��D���53�wjJ���۫*�AhAEɚK��-Pb���Ф��"�������!@DjHLLL\���~I*�(IK�@b �D���iy��^�]:���A�T~UUUN򷻥&;f��+D�u1����qj��/	������"ٳU�@�N�T�vV W���PB����<�;�Trg�����?�3/]���qF���o_�|9I�� Ǟ��@_6-iJ���Mk��;��L"�5��(Oh��m��\9;� �.@�hKx<�Uմ�V\��j����<t�P���\��Gy��#��}kft�+'�������
D-+v���uc�9(�s�,O߇���2����f=G���.0&
��� �����_gń�%�=��D�^�<CήM��t�h)Խ\����G��<H<��������"k0�#��T�޼݁�����x`�̼��E��#=Ӓ����k�Y�6 �@-��ń�j�T�	vw��8%ew�ƹ�dPO���N������K�Ɛ)�mN@�UH`x�����zx�^)���4G_��X1%Ya�	��ۜ��C�L�R�a.7��)�T�����P����u�D*,�|QUQQa��	um�X�?��C�n�z
���z-e����H��P����T��({�z�MW.<��}i�2@�3�-�3c�Ы �Z�"�}��y:/����#��ʊ
���t��мV����������ԫ�F�[�	>=m�R�7�����sL!z�{k`J)�T��p��X �R�����������;���`s�a�E�^�+�]䕽������L����1)g����I���k�j��Ih@'E.�ZZ�Z�+��x���1�.)]9�.���?�LRڨ�OP�HyG�+�w�~C��@ *Gh0��
d{2	�Y�HV���t�N��V�|�^A֪��K��G&����W�̀��|�v��{����44rY7�a(x߉q�~���O�)�?�T2I�����.{TH�S�x����[[�&��XGʯUg<��)b�� *şj�.*�4a?Z��/���ʙ*�������������m�
dP�����p��y>"2�!�ѱ��r�l i�~��y`HEU��6�������]�}��vJp8�������#��3� ZЦMD�&1�NY����d�~k�Q��t�v���U��k!�A��x���nB*rR��xd��
���s"��V��Տp�f�>����D�u�� ������J����67�}�U�e��)gbV�l��(�M/ٖ66g#��C� ��c���x���n���9���ꛌ�>�q��G�vvh/+I$c.����

�}�:C��0;� �n�	��?��m��SKM���y� �[W�׳ �zu&�PX��r���`N"�詩��..��zZဏ$i덅n���ɨx�(Z��x2E�s֚I^�h�&�I;#����ј�Ud/M����͍��)�E�^�F���K�GKS�r.`wKY���Q�z�h{��?ۛ�@&��줜Q�ܖ��D+¯���fg�
�}*SRZ� �"1M	<wK���~v�6�7u������џ}U���СL@_U�iv�/<���j�|Dp�-j<]�>s {(
6@e��)R(�

�*��@�����B���j�,0ߡ��H`y������)(�v\||�:|���R�� �R �6�=ڴ9�y�����'$X�]�j5�	���јN��2]��Ӫ�s*pp=���8
i��H z⛣�iK���?���hV������<8i*
���Ot��ݤ/�	�m��d�FT�7�|#�ٙ�@�`v��Y9�	Í=��oۻrѢ&O�h	\���tM]������NHS�42-9Y��ԅO��C��D"N�єf	K@ ��T��0l�����mq�ͥJ�t�A��	TolG+(���q�`��p�Q��=.	���&� ^.��vJi-��@�����u՜n�K���ъ���J���c��U��q������c���Rv���?��ݸd�M�\Ԣ��vŦ9�⊻�[d2.>��f�׮M��F�ܧ�n津���鎶��v	�s.�*(�*�oo|~Ɔ�	�5�-�U�I�z$M-�<)1 ��W)2VѴn]Yh��4��������u�pÿ�h���	����n��'�	E�)-��{i��m��<9�]�->ƭM�0�@]�򰵷?�Xw7��A�����wT^����A�L@��j�٢��y��6X���{Y�8;���2h9�����	P־>���;�w#T
�"�%遦��xW�S��x6�?�{w2�l�w4�V����H�=JBE����3��S$���S���כ�ii:r�4�*e�&bC��u�"v��U�Ϛ���]coӢ���q�ߝ�)c9p�+:\�?z�YC���z� J��e߼����|��0�v�3)�O�PO#����[Z&p��P�SR�kH��?L�h=�Z�ftr�"�������V��:m"���x<W�a���n�QO�ɹ"/��+)�
j�����PC�s�zfN����f��x&u)��<��	%vo)�������H<�
]��q���ǿq���&Q��l R)���������\��Y��K��)�A(A�}��Q�����ed����B��=��a�� �K�P�m���!j��=���#��_+C�!oB�����If�٠��6֐[UUU]W������T67��m����$��߄�E�qvIU�MO��0h��b�@͡/���:����w0	[�4����~Aql)u��\��_�
hh�H������P�9;kV�b2b�i�%I�m%K�([U1��쫮V����^8�hB�l3�E=��!0���K��A�4�����D!����c�T#���kk;D�Bm:�*g����Q�VI�<U`�ڔnӺ�d+;�aN.��Ɔi�~g���l�'�f�;U"��{�G�);3�i�������E5�.@Y�ZF�!����+>�Ua���\!�����.�t���n�:�#w�`�U[�T�5�J�
���y�0��
y����w���#n��׷�sS���(C��Wa�k
w,��x"Q0C$R������e}��a��t�U��a��0)���r3A=���p� ���������3%���ǽ��r �����
�Hs�f�����j���{V��F��&{}��1+pG�%���)j���i�f󈊛������hhf�'�î(���Kç��j͟�'����D|ᬋu���JjJp,�/Z2�#6�u|��u�>� ����3!B|�s�R���o
���:�4� �ՋG�-*�����ҩ�ɵM�P�Vx�E��=�ǖ5::��������tZGzד�_���f�ץ?\����KEc�3���>���t���~?�@]�gG�% {�ڄL(G�����ͩ�/S�>J��B�P?�(����g����>���*����H ��K5�eZH.TRCI<��?� es�6�T�h=x��O=-`���P�$;���"�ZGh& Vq>:krr�3����4�5%�`��漦�r����E����r%�gX_��Bo>�	�[����utosD ��=r�E�����8��l���O05M�UK�!���� )IH������@\}�Dгo���W�Sk�5DP��̅�&[�8�X������f?�< �x�~�ኴt��t� ��/g����:�䰣�s�O�$��h���BB�fP��� a��s���>�7����9��Ik�J���A�9��Ki0:gڞ� ��)�C�����u�c���/����`�w,ꯆ�އ��a���8|�.C��\{�ਛR|#�Ro�fNP�MZ�?��FYk\�:����p,�=�ʹx����|ؘ��qK�Ԉr�bŮ�(���'���u�o]b_����g�� �8�%�/r0Q+�p���i�����غY�?��\�L���a��������Y�{���o�kE�����.؈��rZ�!#�DV^^��0�$a�7�[���F�d�$ K�;$N:B�R�Vοn���PK   W��X8�w���  ��  /   images/805fb750-7b5b-4a1e-90f5-2022d18e6d35.pngt�eT]ݒ6�qww���=����7���N$xpw���!���s�����������%O�ڟ�eP	A ����*�A���#���'@��,��)F��A\R&�	ܥ��՜,ݽL\-@^^^,6�vnf&�,N�V'�� 9HNRL�;�軗7��@G��#WX���&$2RU=
�(�h�OLR���
	B�X�*�>�z�hP��2���H���;�G/��Ga�������0UD#�� �|y)_k%�E�	n!|�Q�xH��:o�'
�󊳡k���AV��Ehl�atܽ�V�}�-£�z��4*�����R��[C��sN,�4����t�P��P1�s��k�a��[��9Uӳ��$ceoZ���Hd��nD�N���z]`bX��;��n>��v���*/2��Ю+D�Ѕf2g��
ZU#��*�*�Ɏ�$�r\�gq+�R]�P��blz��r"�V�m�BO���N�J�Ӕ1>��Ptǟ��.�;���r84(#!*&S�����C�,�g�"��oá�l�mI�b��k�}�*[�:���rF�չ&�!O1ogX���@*�n��^i���KtW�U�,�p��d��v+�)tpʊ��мb�!�2�L��uh<�V?y�M P��<�	���?Sby�J������Hb��<խ:9�c��Qv|З�͉�c
�:���9�	�(���)HBOT�����p-��b��A�Aa���b��HȣqH�_�ۃ�#J��s�'��L�	B�r6���ul4{��x��i����=8�O�\QF	A�|�&�
>�9�Kv�mb�U��tbDev;ORq�`�o�Y����v�G�P��ˡ���h�3irq2��[�&�����l ��E�lP�骟Mߑ�J��2��E���b�RE��/��m�*�t�jz�Ƞ�*�M�'.a�+F0�6@��.g,S�P�xZ ^rߍ�!*���,�)e�q}	�z�"y�L�bTtE�Bs��$g.������u⾂)c���.ȉ@�F���t�>�b�XC��433�024rQ�I��ʑ��������H���L8�X�o\�8�qgt�w�t��|h7��*�� 	�O���bcP�����?y$S�>���Gb�gT2R��dܕ�u��|F�S`��Gz��)K�jY^��2��Fl������\���o\��8�\G�!�1&h�A�����m�"5��#��
�A��x���+n�<X~&Aڷ�cQ���V!'�졅��rx��}�Elv�4{↽) ����o+~i��K�#\�o�XF#��`�kL����0�TO-�;����"�Ck�������G�f����`b/ ��M��vgC�1|���Ou+�����ܕ�+nR�Q�1�.��7 f ��̫Č_��zE�E7�bc��v�ɑ�*�j	n�g�_&8s�S�J\Y`4`��J����g5%e����5�
D�6'9�eS!�G0���s��s�~�ԗd*@���%	� �[��J���0��)�nV���ݪ4UY$���G��6)���Tư�:�&�X?Ƌ�j����^�bs�7ߺ
J�M�i�S�ZV�:h�+zO�8�֕e�8DlF0�}G�SM.=4)r�1Mw�7��S2��Hb��)UG��>b#
��+0�B��6ϸ�������Y���Q�I��F�b�O��&�Y#
忶�&�A4Պ�@퉲��%�̇���5(b���(����7_�,�r��w[|�6�.$��W["3-��������'27DMbɥGg"yS�&�A(�3`qe�Qѩ�,?��ol
�Mb�KN�P�B��L�V���]Y �@�q"׬���p� �Lg�6gn�::$���/n�(��SʒĴ42��FE}VXD) QJ�|� �7�J&tQ��F>m�wzȥgg"��$�C�5	�:4iF��6/�$r��H{��3p�H�M���T���n^���ռ3 ��'C�h��GT�`�i��m�C
F7�;�V�~_f���BV�?�䪜B9����[�Ҝ������B�t���a܅�oV�ҷqi�t���a؅�%۬��/Z�-����:�B��/�֨�`q�{`9���@��"�k꿚��]�w�����C��0����$F��}�I����·�T��Qs�6M�C1��sX�n��V ��M��Bz�5���&�"\�/}Oto��#�ŋo�x4�3SHI��oWC=�/��@p�r�5�4�{f:�Yᖧ�d"�r4+���({I� | �B �!�{8��;�>��X�@;��Z,��l�qp�.����+����VR&���T�vL�Ц�ۅ���N�<��ٗOt^|g@������s�<�
�K�\�*���VT&�̿��,�F�ㆹ�-�P��4���:��Hy��e�=��f��Y���Vκ�f[j�!�Y<�&�}�R��u�r������V�v�Rݩ�����Ue�Yeu �d�R�{g`���y.�ddd��H��=�s����=q8���^�"l,��R���FJ�@?m��a\��-a*��T*ӛոe�:���:�
p�Z��A�f��T�]Hj�b���T@��1 �ah�i�d"�������3��h����_�|x���o��D�_�Ə��*>KR��뱖CJ�$2��v��fX�4�S}�Q:Q��:pEsR�#c\M�5�2k�̰�CK���������m|+'�dQ���^�(�r";E����;:���E�8j{�4Qsz $M�G�j�@�ä9�ˬ�Y	�׵�w��z�׾���>��h���;�Y'�(ݕ�Q�1gJ���,7f�O��g<C.��$d�� OǋG������Rl���f\m)ts�F��O���s��֥8=�҆�w6 ���]s�6���>�<|h�^��>�R�7.`(��a���gf\�����Rl"�V�D�J��Qh�1�<��֊̰Je��8��1�f��<�mUEH�'W�]er�X�A��hv���N��B9��vWC��i���N�12�X*�f�J���.�����ԩ+��N�cN+��KG#î�t���%��5T�����?�t�$CW�n	(��-�z�L�OѼ.��ƕ1�������(�Q^(}��v��I���(/�-c- 9�?y�]��ha?�R���+3����'�>ﰸ���d���z�a����^=�,�k� AP �W,��:O�7dcrP��8.^j�9>2lh�1�/	x����V
ퟛM�J�����.}񈌓�A"� �0Ɂ�^��U�3z���s������
�7���L������.CF���*�Ġ�Vc�儬vݔsZ��R$�2����`��3� g�)��� 敜�[�����^�3�<AL�J��r�ވG�G�>Ձ�ߴ���l)O�mJҷ,��v� >�z.Fe[$o�s<�F�,�xL��̾����}}��6�q	5����%��1��ŵ�4���=�HB��^%�m�������ԫ��~��ch5�՛�%��YCY펈��X���]�łM�&�"$�,��?�E��.����)��V���4R�\�nӱ�N���l��Nz�h77DȚ�����>9ѫ��߹���F��|�Q���ex!��z*�=
$��_� �y�tʹ�ǈ�Q�L	y�T�sNi�9��Ґ� �yM�7��)O;���)�̲�߽(&'�������W��;f�����=�`A�ivj�=KAͻ5����t���-P�G�:d�f`,��y��Wߞ�U l�x�;Eؗ��`c��(�q�ÕL������Cp5�7��q�E���4�e��F�R��P7�ݚ!U�h�Zz�c�����\���c��?v�cm|��������b^�_�zG��_���5泩�][5��q�J�.VVˣ��A��Q�~F���5��������+�,y/�N;�C1�XSLf/&�&�}��E���V��`��ow6wn��vj��ߚ̳ 8���[O���lԼ_F�%m�[y�U\��K/�u��FXAξ�S�^��xA��F��;��Ki�M�[U��۸#��j�$�mE=ul���Ҏjg�2hɶ�cA�%��eO���ǒg ��Ӂg�����U��մ�*�^U,�3g�{i��b�[����CvR3)��,��r{��i�S��'2�'�Q���R�>��j߻]��
���9((�=7�g�'�¾�V���BJ`^���#�J	-$Xy���	8S�wM��d�0��z�K��}�d+S��}xd�&��mH���@�0.�6�-ǭ��5�1G-,g@��s�boF��g��.����*D��+�A��P:�a�״f.��f���i0�!����J4�BM����JZ��)��?Ի� >f1ev���؜	R��؅l'=JD�6�lFnT��`�oщv#Y"#em�>���ə�*�
��UM_�_�2�pSC�Sx0��*68�]54_��� ��T�V����V���:�>���&L_�Ru��0�,�Ϩb����k�Բ�u�w-���X���Q���l�?T��S�bQ1#.�u�m���@�T����|�9��7v�ޣ2�P	���_X�/�R�j"�O��Q�����A�k�	)i�gR���]
�%?L�{��g���v�x����ZT�!5�%+��ɿ8�Z�~��"E�UW��$ ��+ʊ1�tw�X '�A�=�b�B�Uٌ���xl.a������|0	���	��G/S"kCax@��8�*�c���C|��	�z��7�7����� .�M����׽/w.�}�$���U�y)��>��US�PV�js��qe�dy��yo��<���L��F��E��|Yj<Z�b�z���0o*��O�Ƀ�4P;�v)�֒r��FTIw��y#�s2�6�N���"c��]ψy#ɟ���b���٢/"�l���۸����IS�0����a:?��B&)bl�M�<��pT?G=)Z���#����Ŷ��4ۍ�l;tXW~L�/7��볝�ϩ��t��_�"c; �������«�_~�_#�k��&+���>Be+�o�!mX�rX���x��hޔu)���2�B��H�ĭ�g�uë����j`��R�X+m��צ[�ւVǫ��:<�p���gtU_�(䋎��pP����}nMIj��?��L�A��n�?85�2�?�#��WQ1:��C&1�28j$�{tx�%&��\�8fvW�<�)$�S����:������?��S�h��#mx%�s���W��9�K�w�j���m�*�� J2R��vx!��!]���#敗�緵�Ƿ�����}W��o�!�#�x��/$�eX�-{H"�UܯAJh���<��hEq��;��OA~�]��0��ĢB'$9��j1��h}d��8���3���šg�:�c��W��[�A�$����}��]�����d��_?��"�o��O�y[�C�0�������Q���+�^ppMu`��7� hH��������������+����J�ץ!����M��'��H��S��?Kϐǻ���gI�1�kՋ���B�b�u�8�4R݈q����#HM75��Z���M7w��F�5���͌Q��^r��׫	�m�v�i���93�Ot���_��.��ٟ��.����8W��[�ǘ��(W�Df
��R�Ո�gL"C��v+�Iv���Ý�x"�{H;��l��9����R���`��ߩ�N��y|o^��ؓ�EҪ:�+�#��ɶ�
��*�K��Q;��8�1x��YU��B^¹���yR�a�BA��/o9��MqxW���>�@}:T	E��M��n�&��V:���g�_l�|0Q��m*�n�&���2���mSeR�&�cx�z����	���6�Tx�S��i��=���?������O
�bc��0�\8���L�"�ˋ�n3���t�O�,H�e�H@~W}͏��P��V�+�T`xr)�TOLb����T\���1 HWQ��ʃ}��ԫ�ŝx�1����y?|'x��.���٨�+�P���z1.�����>*L�,쯅�$~��"]O��N$���p��u����"NF5{�Q�m�O������MI����j�d>�u$9��|g� �h	�}����,-�\m���\ѦqV���M����/���7n'J)��Ts�w!�S�5��aE���\Yr��*�<�'O11�Pc&��ߜ�
K����Ǝ~��NB������Q�����@uf[߿�W.�`���Z�⤀�L$:����m��O���|o��{Ԣ�""8ȃi�M���á���wm������c����䚩��;�tr�e�Į��T�q���6I'� �4�u����2 W�rY rSin�����_9E0���4J���	v�'\5��N�ˠ�*�3(�� �Tߵq7F����B�'^-��3��������ej��RSv� ��>���o�M#1���|#.xmon��0=�3F��:�PE&��^BM~�������T7�&�fWr/9/�1�m������e�`YK� �.�k���0��]�+�#0a��V2�ZBh����#�cO��U���#!N�`¨�Tu������]Sܽ��K]Y��#�7�?N$��?����W�IT&Ҡ��63�j�yn)���$}�><熶u�ߚ���T��.���;7!U�
c90\��mx�.IM-�g��k1��w�v��7e�[��TL:�����!�+:��i3���8`�f��M&�VH 3�[�d��$}̯�"�, ��#w�ϔ�?�bcqo�)�QL�6�2��3���jԂ?�vk�i֦��ja�IM��qb������(�$P�N���Ŧ�J�w��M5�-p����?�Wd�C�o*����ȝ%��3�TjJ��f|5�m��,�T�w+X|x� W7���*�C����N.�8
T4��}�T��	����6�+yg����f�z��T�/���*F-zj��&sU��/��3I,/��)v!�|�ĺ�t�=�47�bj����k��4wv�H[9<�1�ރm/<�R`���T`S��c����b�3�����L��4�	5-��D��� �e�w+z=��	�N%!���N����j��%�r��O>N���8?�)��I,?3�d����K��j��J#�<4�b�h���L~��S
��\��v��
-/<=`4��i��7<l�*ڨ"R�,�r�UFU���n#Ü���k��;�D<��A�����j��} e\@��Ж�R�����Sh�lzU ��t�jv�ۓS&'�V���d.�	0��ߋ�o���}�H�c��ešA���i�U�����C?O'�ԑ�Lp������r+�P��5b3��g��zz���5~b���`���q���I9q�}
l��J0�L�r]E�1�c��᪓��?�=��o�OzU��s£�NG�v1\D"6E:���a�^X����D5hU��W��L��s�DV`�0�r��-p�g1�H{�@��]t���T�� 2U����5(gd@����K�*iL\}G�"����pQ�2l��+}&�Z���9lݠ���ʑD�|�Uҁ��[bed��Q��Y{ű<O �FU�:��	�?���c?��T��*�h�,I�@$7�'�eɪ�$�XL5H�����2	h�8��?n����o���Lf(�o��0�i�8�pK�^�����ȑ��sa$�B�;�?s�*A⃗�,����ݓV@څ[�(�!��wJ��|ğ����3���o�6Y�e��&���cp}��~�#����?ҵ�"�&�*��fETО}��tխ�Dq�Se!=��M2[ĉ�����k��]��y��64�Y뱱�p����������3��A��f&�\�$J�YOW_]��#��ʏ�t�)�s��3}�-��eHM�]�?�-��fkOn�M�J09���J�i9*���Y%�"��䵂ڙ�w��@wf�A|��x����j�H�rn�j[*�q�l���#jzS�B_��U���T,w��`�OM�ٻN��pC�C���	I:�*�,b���:Y� �C��<��PQV�=a��|'�<�B��.e�����a%�i��2w��]o���>�{�S��u�3�1�Nc���){��把g7�p���̑�	�B������Kc�����2�ʵ��v��[��'vz�#Ó���}8DÚ�k�z�1�ᰐ����Yko#nc��L���I���%�����h�v�B,5X���%���T:Ɗ���H�u�����p������!��r%H��c}�x`s�h|���ߓ��\*ɰ���Jl+��c�@
�|�z��f���-�&��]�i[L�!���`	���q�yrb��㘰�Q�C::����r���l*�!%geЧ5�f��O�=�;�mC�ެ����S_M�J2�����(�k�#�Ō���t�3�%��e�WG��
<�W��_U�s������c�k�.�)��'m���n`0��U���i`���/Nmp{?��g��no�t��\� Ǩ�F0����x�B8�O�B7;!&Nx3���1��
��>�U7�R�K�����R5��w��~>�%_��`�G���(z�m/-��pC@%��ij�H����$�E��OFH4Xj�J���A$���k~$�e�}&|3.�G��ʺ5?d_�{��z� �<����z$�\-�si)s�`v6_C�p���]^-8��h��yzv��{�[e��aq}���:�wvgW��m~�?l�do���ZN�]�ϝ/}�x�����ڵdM�m%�H:�7ܵq)h�MVk�>�{��t꽼�\"s.(%WLjU�j�֥VW�e@�K�9ޙ}��'�	f�|���-����͍���(�Z�s(�r�ӼA�D�����56v��9Ͻ�YMڈ�-@h��=�(K��$|!����]ܗ�ά����n&Ґ�`�I��~R��I3�ý�j�'^N��,��E���ƞ�I(����	"��� ??�����v8	-81�/�̎M�sj�,p�.���d���O��亜�D8f�����fM� O,�� �GAUϓ���4�2�0:���b�`�q��]O���]�Y��`� �E8�{��S��Yy5��l��e�)Q�I�։���3��+�b�{�����3��fx`lltY/�A���������zW�w~�Y=hn:��፛?�b~d<��:��S��u3U�m�U��G���������A��h�� +�~��*�F��4 ����J5'!������ta������yn�
e
�0��62�W?t�oQ.ѱV@Vn,?*+�c	�s��T)i	�����"P �{�-ݜ�c5e��F��{Z��mﻡ���
���ۀ L;L:O���}b���oa���{j�ߝ� ����dtB���eѼn7��pM�5�����{���Hd���l(��`�A��LBQMD�F|�iw���i��-�b]��͂��p��P�nY@���cT_�.Ywo�������jID�bh�y�Q((��}����h���}��� !Gۈ@�ȁV���C�p�0πɽմ��j��{�[�Ht�m4oJ lŘ�Ǽ�T�?�*^[de%y>ɐdS;&�'M�����t �W/ט~R�~�k��%�؛̓BDT�l{U�<�[��%�����i_ߩl
��B��E����zi8=kY�v��$�K���|ۙ#2���dɳ��i����@���;��� [L3À
��&��ۆt��5%�e����c�~ N<T�9y�Vo=+X��Ei���g#���\�d�9��Čp3�ݦp}e�3��>}Zy�N��z2f�m�c�~��aF�>KȌ��;�Κ�̘ؼ����c`H�ҙ8d��	������e����x�#�l�C`6�Ҟ���mWge���Z�CPu>ts���R�%��Ȧc��]�W��==��k��0X[=׮ߓ��N�|��+�^b ���o�Z_G)�3W��j�92�l{(詭��y:����n<���&{M��acpxHBE� �P*�&�����gO����q�%9D�Σ��
^:�1���,e?���LwCM][��iwD�v1<r53�$u>��BU�ҿ��_'�$\�R5�9�v5�7;}w;�m {���[���G{��nD��-���l�^6�:nj��ã��7�=��[�݈��ib�IERCٱJO�&�۩�.�4�-H&?��7RK�-����w�Ԓ�c�����(B��̯"��
�������Aۙ�0��먝���gdЊo�	�˪��U����z�·����c� �_\�k���c�-�2VpC��e
zo0�����1Ds����s^��Og:��f�h/�[��xU6���#���޼��ɞD�-'/H�\��a�l���}I� �G&�j�t�sK��g�bW��\#�=�� ei�΍��4���� Ʋ����VI(����u�f.	����I�����k}���ʅ��-�v�:��I�Ѯ����<����x�=�鰘#�����l���6�js���T�i�N"��W{��j�h��+�ox��̻ C���)ѓs�E�pzx�͝]��q��J��͙��{j�a���j��+��l"��΄.��+�[��9��s�*����P���]��z�s���fu�t��'�ZY�5��/4m>��$�.ӎ��`���{'�ǋY~V�R؛�(��O&}��g����N���ڐ/6�v=f��(9Tl�rXQ��� }B>�9�6b�sd@%��� B���y2W=�.^�^Þb&�^ԫ���Y��ؗ"�h�ܪf7�I����d��l֕��t���?�3��8S�����Y�󭆊��x�^pNJ����1��Yǂ���1�:s~�������@�����h�a�b��%�zh�a2��hOzfl���G�e��ӟ�e&�58��Z� R%v����-���$�O�_T��s�M�e�>�{���{��Q�7��h�9 �>..*✕=�[j&d�7bz\x��P��r$�Y������Ck�7ڌ��>uK��d��|�6�ǯ���������q��L����9Z����q�j[��6�.BZ6�_��\�� 0�콳6�������;�|�J������}y̞ޜ���ޟ����t
����Vj��'a�׈�BW����=�@|k9�4�W�G�,q��n��~ӺM@���~}v�EY�΁@�U����B��ŭ�AY��―��=�Ps}��V�m�E�3�����H@�����S~~˄�4��|u�խ��-�����Q7�L�fTE\�|9������� �*˻N�@�)��
�|�+˔��x���P�M���\��������6Na;���ĵ@$b���d��q�7n}��1�^���cBW�y�=�_�^絶����*���q������� ��ǣ�]x�� �҉��Z�>kN����2V��%z��d�t�󅹌���Y�ـd��<؍//�Z���A���v;�>-fUy���yz+��ܾo��sK3*���/�&Z<6�S4:�s�U�V;�����<�J(&MF�'_��n�&׋�ʭ@��?i6�������nk 2�֤�b3�>��
\P�\�=~������>�DG;X���O{E>_ �
�UV��@j�m�A�����p7-�������GY�q��^
���?�n/�\Q��Y���ڒ���|i�"C����/� k�C�6" 
���9�N򕡕	�8��IZ�x�iO��G��0gD���
@ț��޷@����^h����B�o���v����S&����!h�]�" �4i ,[ϐ�����{Y�qc�&[BA�2X��8�x{�!<H�'�zά�G
 4�;�r����� 5ҷϘ�4��j<y$�ueB�w��P�ԍ�p!&���ߓ�<Jb��^��R�ޏ'l��P��h�-'-�)�8]M �L4���ͬ
��?u�b+��q���o�̑-nAy�K#5S�a,�ˁD���鱃7Y��[�=��Lޯ��ָ��h���L����ۑ&q�}�[݄ɞ�Qvv<T��n^��&JF|�r����H�����Wr�;�h|��"}EH"r&�0H4�L~\����
��.�E,��v�_<��9�B�Q�8����J_~%�P�n�h��l��e�����gN�,ը�
�����.��w�����5&s~��P�P1{�7^�D�v�����P)����C$�������:R�6z5$<��!�~$�����h���[S��y���Upm�JI\��k�6�f��A�Ɵ���vF<�?��;�q7L�]�M�1��b�R������ŝk��V3���WR/旘��Ɍ`�jQ��J:�t�$A��[�8�=��<����Dc�z4:���O�P���t�/�>�.�ߜJ�ޕ�:��1�d
�i�a�,�����3�7�8jH{�,��.��=�v�GY�-{�ޏ���~n��5��ΠMN �4��z1=o���m�ZG�.�l�An�[������`�!v��� t�0P޶y������{|;n�
v�E~#�����-���4��[�?IO\�X��t��S�����\p��oHa�t5�b-Էd�u��U�:"�4�>�t0'�Glǭp����<���r-�چ�p4}�<a!��a�|yFu|��K��N��z�  ��n����>:Z�ĥ���b�M9����BL�\�������#�~ �i]���]8�ݏ�:r{��y�eN`f3{#ާ+���k!����U&�Lа}Z·:�5?Q0HqÞ#ޗ�o!�]FU��8�5��w�TqKq_}�	c	I�|R�D��&��_�l৕/���Om��w;d��0�wfKb�����y�(�(u��\��u���Fa�������L�A�\�_��jP�bPihX����k�!��I�y�eA�9�f[j�3%�_����M�T?u�>��ru���c}/:Bz��Q��υ3��=�4�d�g��0&��?�>m���FȌ2[b���6��6`���(����^8��#���l������۬��&__d�s��_��ӎ�٘*���oI��8M��,����i$�5#�#�� �c��,��|A����2Oӟ�&�'�6��,s���z�����/;�G���.�Y-d�}VHYݍ�Pg�Id+q�Q
�}���3��J2��F:弜�z;�yVU��������.g>�u���@�;r���L����,�ɣ�DԏM�Z;��F��J�IXb���cS��ɍ7�*�RX������+�X��Y�_��a����������|xg��q�7�u�c�~C�eY����C
�]@҄7��p�5�4���]}��lɑ��
yv�\GG?��fz~��*�Ts��x�
���u�]�k�W��Fч�	�Q�������W��׷h+��M�hftK�3<���S����7��|!��~�y����bIc� �v�w��cb�����S�J������Q�������X�Сň��XI��퇇$�߼H���~� P(u��q�������T�L����9�dm�ë|fUr:Q�QX+d�^d$���B����QX)�q�G�+rrr�J��x��u/�}[��!iD���[���KQmt"�Xͣ|��5��]���~�^nc�u��l��c0J�o<�C�����E�k~	�o0嚱{E�>�L�Dp*:j0��_LE>�Fq�o�S��fKگV��ގ��yk����銀޷d,' ���!�
m�37�^�4�1��8;��]rfd�:̌X2�bo	u�H����E�C ����&�2�2�W�uE�J]��\i)I�av�|=#�Z���ݬF���1��Vxh8��{�l������ޘ���������p�����f��_�l�� ���znl���A��C�2&�V���7+��!����f���9\��M{����-����>D�"��[=Ku�@5�i�H���7�8L����:�۶0���/.��3:���fޓ�T�D��b�e��[���~\��S����%@�����͔!"����G%����$z�)bw&�v��'ۆ��7�i	�M�T���"����c��jD������LF�F��
�!�4�[t���͐�wFd�o�T6��s���~���f�Q�I�s�����M�
L	i�G�Gٿ�T��'��ʴ��~r��ƟLw\�)����\uN�@���G���M�s���	�̥�M������[M	]\Y��U��d�2�a��$qv�� �<ǁݑ��
hV�o��(H#^X�@T�d��kl��ZW\G���\�D���Q�>6
Ѣe|ǈ�R|Ȃiߓ�_�Y]>�h/��I.��ՙ>�p�g%�-�5 ����g_���&Uӿ�4�(�zs�A؄���ɉ�Vpj�E1���x3�p%1����鈯��vBʅ��F&U(\w��|6a��IhDI|��[�1Z��D��i��q��}]��ߝ,�T�y���ݾy�*�7�*��n�F@�������<���ε�*�22��$~��T��h�s�&]E�Vo(������{}��
��o_H��.O�] k����DhF?�n�YRq8�(vn����0?����`��ƅ�"o�̥��cx���E�Z]���l����@.dd�)M�c���D�L�k/�\�>"Qa��K?6|��q����ff�i�y��XC���Ijq���>�Sg~��hr����ř�N�f٫	ܛ�ݲ��~�1�#��p$�yؾȵ�s�����d5q�=�,���t���iyN��Nj��tL�/�ﶵ���ɉ�e'�����vn�,�·�_Y��s|���~���t���{n0�c�����ŢR:����݂w<L��*�i��\��t~'�>Y��f�aPꔴ^*Uk!��|4�����@�v��A?G
h �����ͣ51���/x�3�I��h�_����7�*V+t��]����F�v�:OLM�}e�$�����Fv.�͒�O�R�<���u�F��㖩��?���h�6.��"���vkR��5�JYhh�5E�W�6Z^���[��)�	�_~���3CB=��9�(5���������� ]<g���������v��8U˕�Ӵ��{�nӺ��o}���
�o5��a���� 2�]�E���5P��cl�n���S�6_!V�}�#��bi�j�h��Vԋ�Qo��8�0㓲��._n���7��aD����C��1���ɱfM7n��k��;].j�k���#2 4q��7ȃ�̝2gM���%�G}3o�C&³j���b����I�Jb�MkZ�i ~ g�>e(�����������ҙ�7/C�Yd�~Z(5�7Ii醆D�*�A����]��X%9�E�Q���w�[�q�WST�A%+�-��/t�b��I��������^�8��X���L�{���EX����`�>�1Y��$���? 8�M��gP�����{�#���"/h���NYn����7�W�$hu�z�KN�B��N��� Ѐ��,l���f�b����gkV��5ӟ4���O�pG��ø��s#�����>����.w|��Q�LBR7:���O�Mݽ)]o������k���s"�ΰ|1:��f2O^�����H4u�zGN_���p�����Z�^�?�x�b��������v��`�<�h]$�89��o����sf�
��2|�S�zE�����e$/p���`��g	�s�0R�ĳ�{q��Ӡ���,NA�����ޯ֓e.uǹ��*����{���_K���qG	�2���eT#��|��Q��N� �3��C�Ņ����[S���hi*��8��L�
e��R���T����sV��3����j�$m�`g�Veۺ��v�R?�<����C[�5x%���`ۊ�pq���"ph����in�/'�t����{0>�����AZ�V���L� d+�4eO��lԨ#��^"��܏�ZK�7�G4�����.5x�Ά5��b}ꁋE��`ShQgͨ���-j�&��v�`VC�+���J��z��9���"�� h��F��Ӷ��D)亢�3�q�$<݀�5D�x!"w
>��+�.�H;�h��/�����{oCۺ-U�縯�q]XX��Rk ����k�ފ�������D �`���.�x����m�%��x	��>�["���y�ǲ��LW*�I4���I��!��)f�� ��G�m@ze	��(ح)��tX��n�cNy��Ǎ4]�?��sH��E �#V��t�Jr��z�/b	b��c�B��;��w���$s=�~s��*U��Sc�����!i�5�����2�;���^.ߏP�Nz�yE��ゞ��=[�9$��y+�y>}7,�mw@^ͼg�����~{����������>xT�ݺ��#15��1�߃K$cv�"�q��O���zn�~�������v�/b}�3H{��]�N%�{5�}������4'ec�L�H+�8�����!u*���)��_�NM6[`!-c�FW_ 
>wH�n>��Xƴ�j��3A&<��CI�G����7 
��D�+:��~�p� �=���,���={��[����0�%N�|���Jj�O< �I�\'V<r��(�p�z���&~��S�e��N���*�xo�*�ǉ�wg5� {�ۏ�'�|�d�.�sc�q�Ƿl�����j���EAT�D���R�w��+H�5� *ED@A@z�%�BT��tBh��Jh���A�s�c�W�=��R�^k�������=�,��jG�Sen��S �ۻ,�K��3�N��|N�!|,�|$�ΜcB�褎wI�7�i�$E/(	��q���������U/����l��mM�˕i���r�)�H!����]ߡ,�-R�P�{�{��{��k�ec�d�4:���Z�~��?����G� �0�Re���d�
߬�SE�#��G��L�X�W��3y��Nڒ^�P&؞y��/D�L]W��ȣn�>H֦���aF񎩯/qB�	h�:�?K���U�O�g���.�nkH�����³�;*�2�3��a�!��G�`8e�5�)�-��q�������u#
��I��`�y�:����t�)Q!��S��N���k�5Ғ=Y]%>r�F����=�q�\��l��h Z����% ��@�I�]���!����	��"���!�6�@ڵ��@w���7�_�C:�M�&��-KFPf�1��!�n� =�A�ۋ�ҋ��Wyy��ӛ�p����5��I��8 ����!�D�����[Op������\���S��P��@���k_zE��I�n~�1]��lI*L~� ���R������BZ�x���p��>v�&�����ʒ���R��K��-�~�D�b�� '�<9��?��E��:'�o�����}��H�N�C�>}{J�F�iL��9��  p�Z�G���^m�J6�ӏ�e����؊�zb�4_�2������G*�.s�����}��0إ@�$��;����*ʎ<&d�g����[Q �lK��'^b�Wb�h�n0]�<�����e4���O{�:�^���I�J��5X�M@�GV��}��G��c����Z�����ѝ�N��BZ����B�	�|�R(q+z+��F+}ނ�M�jaQ�d��U�|^��g?���6��z��Y���מ�M��<�� 1h[��xu����e`����)BH�$��٘F�r1n���)/�=�qu%XC�+^2߭�R��v3K�1Cu>�=��J;Mͻ��Q����ܹ=��)Q�\�!v���SE�ξ#�gs����R�T�k��}-�i�3_�n7��)T��B�2���=N�뒼���Pza]v�m��ۛx%������/�o_�Rpd��X�ʞs{��@B��ok���N�:�J�}����Cx&�|��5J�qN�) 4�P�W�����[@��(�>WD(jd��.�)t$���Y��T��3�)%|��b������
�>MFq�=U�>~wŤ���1�\AZ(B���_�O
��x����ܰ�i�WPT��n�s�ܴ��#n�Q����!�n��۩xܔ�%�gT��Ǘ��s���H-ҫ�Tgʲ>.O����Q�a���VC=x�{�T�5�jc\��ٍ��X�-
��-[N�6x�ΕbeHvs����A��8-���	e�k����f	����\cD���P�*�:�=.fT�޺k!m�
�F��-l}�W��~��	���Y��#[�ߏ<b���ŉ/	�Emmԛ��&���ў��eԨ|��)�r�_�A��b�a�-RSkH(�	�GB�cas1�A;���U~�0���utr?�\^lK'�`C��wi�\�&���{�dAc��*S?�9����f�w��,J����^>:��,l!�8yC��<w=������))3zњ��:�l�s��:0��ycm��cB�5|����<���7k���b�ל؂�.RK}�?}�]V�����kr�����9��}���d�TT0\��x5�k�g��c2I�ӽۋKK��gU?������\Ն������*�Ŏ^��r$�zq
7vt�UyoF#�RR�wM����I����{��A�C���h��a�J�[��":e�����=8���T���?8��2%���������'r�ˋf�BZ3��BZY�h}�|
��&8�>S�.�o�ͻ���O��'������m}5�c�;X3���m�zb��9J��2R��o�����|% d�xq���_^��y������{��^�'ĿxBxI�⛇2���H�L/>���#y�����jh�~���%�z�i��$�j+�'�פi��c����N�io2j��yCM�y�)&A��|�U���U�~RH�cF�����=$U��A�����$	�����!�ǏWu5�_D�{��F��Ab�8�t����1�1�]�������s�2N����J&�B����'��4-e�*~~�וh4dF�k8SV�֖.oe��~$���v$T��O�/�R��뵠��gМ�:t�JE�Kŏ�c=�&E��i�LaZJJ�������~~Mj�"Y�)Bʱk#%�D$�?+���PX	"I���O��L���&��&�˙6V���1�k���_RR������������G?����=9�cb���ϰ�������y`���ڴL�~�q���}��Xf\mԸ�Sk�����  ���`z積1�=i��^��,,}�Si\�OĬ%RhR�t0�������w$���6J��PEͧ����'����V������X�ii���҇z�'��nP\����*�����3�����Cf�����9�S����k�����;݂�P-���4��O�'8R���Ƿtgc��ua~s�zo�^�ώ���djr%���au�gm�O�jZx`�^�˼����^��n�TD%Eȱp����g��(ی	+/���܄�h�m}��<�J�K����0�d�{L^vo��|؃�6d6�F��ϣ�����N=��ᾒ�;�F�$'����*�ǹ�a�G�5*
� �&�^i�Y���;9�>����4� �t������U	�G���/J��P���b�?��΍'�^�lPT���xM'{�?�ka����%�{.S�'[E��Z��ۛ�cy+L��ʵ�2��y�Q��ڇI�ݶzm���B��Q�Mo�X��՞�Rl����%竤b��;����0�%���	���;�̝�Ȗ~�e&���/���L|�^h'��ш�q�y�3|�1�  iX�z��\; L1 �e�̩ķ���71��qx��C&��_�,��wML����'���k?��ܨ�zb��J�C�p�C�|��#��>�8o�l�d��P�YF��wMsҞ=��h4!є�bY��棯�^X2�'m���a��dK�n�NJկO��t��ĝ�QKL��t���+��#�����"�7��\�L��%�� ��J=d��	�޽�@����Dp��14��B�>����_"�DMnWҋ�*���@���k��N&#�ʈ[�ѿxp>]��f2�)���DY}e�3��2)zQ��x"Ϟ����&@>խ^*�]L�TPX�ſ���~�w��łR�Wo���'�v�%�=�)b�׬ H���8����Q��j�"�;
�a]���nP\bb�EL��:WȲ\6Xy�f�T�"c���{�/
���������g�=b-YZ��ؓUX.��>��T��U:!��x�f9���DHL��6��)����Ʈ�:"����F.%jp�IG�d��R�&����a\z%�~e�u-�!����)�7�Xa�JGW$����e�P��&�FGǎ^��,+�R*$��Fo� �~�	f��J���<~�M�vd{E�իW�7���Ĝ�솬w���D\�1$T�	�L?~��)J�F{�1~��O�Z+T��j&�@yR��ro�G��臥�J�d
�j�ڗ��L�NTք���0 |�Z��H>���=P�"-����\*�U�k����;����N*6�P]d��ؙ�c�Qd�`�9;� �[�Q�֐u��S��O;%N�5�B�+[��Qʤ�� ��}\�yU�����s����Z�ms���cx���"g��3
O��t8'����@x���
y5��v��g2��Z��s�A�+z=��`�6�Jۮ(������I~��%H����>�/u(��Ih��ܴ)���>E���r��7�f�7�M4��3D4%�����5���)錬�L��?*���u-��q�"/�oF�v�<ο���\���Ԩ{8�E�����)&��*K;�����@�l�)���_�6��܌p?���.�H��0�}o_�'�������Pɋ�����j}$,ژ��_����n���G.Zݽ�&�s^X�ouР��855U9jy~=�F�yV�b��z��տ���zl�a����1k�[��k�ɩq\��U��߼�R�9?��df%�����5��uf�իWB�➞�x���#<k8���8e%%=�0����p4Z�:�B{�5?l���$'�[�&j��;��!i?��^���H$M��p	����A*T�â҈Q�mT�z|��GpW��L%����N�y'��͚'Tu���oJo��)�=:�C���Lׇ���M���,>4����~!����٨r@�@����|��}��?3=r�����/�����dYe�|�ʓ��C�O��	��������Ǡ����6�vj��㗷�5�{��Ւ؋�I-#L2A�ɡyMPr�gFщ��Pr���ʶ�ӂ�d��������?�N�!W��""��x�O �^&���|�v�J<�u�l�r��F9C��#����g|�M�۵�#�:��M����/���|d�����LÌ�|o�krW�w���z��>�:\����Nx;�TV�8�@<~�,�y|o?v�GF��������U����'�ċ]�Q���>3� 3���7�@�o��̟���D��Eb��ŕ7g��>D���@@P��X����E��`�V����ʛ6������63����C�7�cf@C�jt2՝#p��X ��x7ٳ~c7��1��W?��r16ˆ���3o�?�m�ZKL��*�����U��{ITm1b+����k���]|���Sp�� ��~�9�ؾ\�׌g0�������;�%����	g�UE��f�X��7��}�k`8��z%��ǧ�����r�rm���ݹ�oy��/�V+8�G�F}-7�0��~�;� ߯�V|a��4�+�z����X��M�'�c d|��[8�M�/��2�� Zெ���RN���Cq�!�/�<=Q4���.d�qOqv��+�>�_���>��R>�D~�$���1�GE,h��MP�����O��wl1���Z�3�i�� � f������V����y�?z�Z�U��\h��т�r�f7e�������u���q�[�5���O	W^^��a-�X�V�A*?�^q$.&F�3n�Vl-����d���#Q6�N��1�he�g�7�ǅQO�q���NЀ8��Y�;���69�n��z�ZQ>���!́G:^/���5�J�~nz��H|f3�mw޴��dSP|zc���KZ��m/����V����C��Z��A�b@@3	e���7"NɎ�J�˅��5�:�f_��߹Ɲ��5�w|��Jf�bW'Y�9ب�'�εz'����PΏ�z�d��74YM�*�:�܋�GG��"��+��mx2{��P�\̤�&H�4�"KS=�Ye�;�CIE6��ƴ���ҵ(D��C��H��JM+�e��:��+xݦX��9OL����"-f��@gBO?P�$����o0��"���������u���-)��wPi�ym�OТ���E%�Oa�p`A8>��	A�	~��7��P(�N�W�A�z�71�=��`6X�w2�f�BO��*	���Ϩֻ���]y#%.� ���VH�g��>,�|,V�uU� �[���P�_�eL�_��Cv^�h>�&z+��C#o)&�\[:o�3�6յ[XR����7:�5�=�ES��'�?[��`�Y���ܻ/����������g6 �52zL���^[��i�SW _�ݞ�O<���32?�8�p�&��D�&�щ�|j�scrv{@������QL���y�@Cu��G����ϿJ�/���o�)o�Y����>r����d���9�1�>�v��� j�����'�1�I��B3��Z;�?��@���m\�>����~J���%S1$���H3O���Z���#r�j��5*
��� w����V�.@�m����HVO����s�'�x��y{���=^r��Gj�U�G�"��}��Vv_I
�B��T�iv�����V�kQ��l�?E��i�[��QM0"�����1��̬�{3ѧ�\OaI�dl�$J�0��k���'B�a�' 4��))�)���]�X�)��w�߲��ON�|�@��?��Ly8C$IM�T�c1x|�3 �K5Q/[��N�����{��<v�%�uq�]]�o�܀���++�q�~$\~#!)����cO���홠�m)ҧҝWؿf�"B��6k��P��րχ�1��Wi͟�o]����-� ^ׂ=HT�2���^Ȗ�U������˼��ݰ�-.|l�=/�(59z�oJ���pY�ބ��������o]�(ص'3��ֺ����}�IB�RJ�Ѣ���52`zhH�TL�H��~�A�d��4�+t��+ی	XմT���B���[��\���cn�+u��mqwW��R���.��M�zg��4� �E��'�����l��Mtm~P�G�+����v���L��=�a}[����	SN���c�/��#�ӊ�y9����[-^�'�B�c�rNVc����xM[��%��!���.�7��3S���ӥtr	�����&#��=>VK\%���T����ƞ�w���W핖�E���P`�zHUȗ��!qK�C�(f7�Х߮+���9�a{?�B.��Т�@ѐ����U�2����uv*n�T���gJ��)��,�Σ�3,׸�2��;�ds�V�_>����`J�������w�7�j�e���>,�z�����+���N��4�(�z��I]f�S ������r�ʽ	쉶�i��]�i�댲�����rϙo�=�m�e�&#h���|�|�$�B}u&K�� ��٧B�뽖��'9u���ڕ#��s��r���]ɓ�����>"j�NQQS���Ŗ'K�V澷���tI�kv|�(>C������%$'��Sꞡ����J󐇛�z�N�	Ʊ�<K�ڼs����3N�'v������ַ����^�Y i�����H�`�����G�b�k:�:��}����\�"@�]�z�iM1�mH4��3�!��,k�Ԉ����b�_ִ��+�<7?�XCtޤ�ω0�5.��l"x�F��C�C���Lm�X̢���2w�8���i��^��>֬a6z-b�R8��d�gZ��Z��z���Q�jH��5���v8镳2ښj��֋RR�M����ץ��J�yp¶�{֮�^�b �.���7 ���O=�t����D��F��5b0G�$���y|�ܠ.-��U}����Y�[¨G��Y�bHz��K��f?M5�Y\��K��f'�������j�q p��C��H��v��K��j�6�Q��C�f��qP��Sm�d,�.�:ʘXs�F ���;�ؒ��ҽt��L�����)�M���6[��h�ëۿ���,\��c_��l.<�?�N�<��̃Tb�1�ǒ����ɂ�q1/���J䱇��tͻ�{�>c��Xr�X$˝ӌo7/on	�7[�� ߫����x��8�@��ZѷOƸ'�l7��`vR��G�P�5@f@��2�D�'6��X0�m�"O���R=Ǿe��R>:i�5�|\�r�%C���LY���y����m�-S[�V^e�*s-���_�j�f�Dآ8{B�˶���T��ĪϷZZO��k����]��M��*��� �wl��nc����5�JO������$����6�(�M+z�҂V�";���Ϡ��W�p/�d�?/�R
��ʿ��^�pH��+��*���5zd6K�	��iRe8�$l�Y�pD�O��"p#�|��CA����#T��1�C�)V��(1��Z7�upߙe��Ρ
Ł��1�o�shP����p�Gkmkjzm�z�����6��V�������5��:�3��j0���G!�1�����Ă����>�����V��������BN���K�C9�F�CS��j'�YD�����=U��z�*�o��f���.�[B�9L�~�#7�#���:�ܽu��Sr)���go���w���h�v�V�)xsʿfr�P���u�#O��v��5(��G�4~[ЪK�҄�T��xu�E�wWM��|6�R fs��)"�E�c�֏���_�Y[/�4&�|)ryef�޴��L�=d�`��A��=X�b�M6�W'>�n�>j64���P��@}�L��&��!�%t���
�}�����_C�Nq��q]G�T�G���{f��l	�b"��jc�Z籟�R'6��&|���>)*�zJ=��p/Ȩ�7���fKve���L�"�r������<.�Z{��ؑ�IR���A���>l��������6�% �r'����6�F�Lw�gm��<8=SQT�ez��\���QY���u/�Y�>;^��\Y��<�Vd^������4��*@�<u�4�[��	��U�1Z�pĺ��b�N)2uXF�]3e��Hm��=(��V/�f�n-ߔ��������n��6��:�r:����]ss�ޯ�o\m�'"OM{{�U��#����~!���t��%#�>�&�涘 �"��%�ٞ�������IZW�o@�_���XԹ�x� �1	�׹�ܼ��!���N; �*��A�>�j�B�<�9zۦ����+ut�>ɘ
۽o�-��q�����*�Dŷ�b��@+��)��K��y�[�/GQ׈WRS���x#�Ej��Z��㏻�����r��]Ex"#�"*�S�N�-�Ddk��g�#j�Ï��P���s���\�-���˴'ּ��tЇk/0���6�U��eA��>�s���?�9*�ϡ���;rh�.jz�{n���,�#�|��l�c5	A�o�
������67���e������7�p�	Uz�2;��I���,Y�=\WO�YEc�ײ�ȥ�C'4��X(��f��k�dT�E)��:r�i�nX�V��^�s�Q�����Hl=q�wz=Qk�t�
�z�P>�EA���:+�U��a�о�}��ﰠ���-�@$�����\��<9��%�$�s
��+���P��,�R�ʝ2\��0�}�J�f��Ipꨣ7��x�@�؉Y�������g�o߰��ի�S��hV��Y��=bZ�{�i�t�&F�K�/�u���t�3&��\b����V���W�fN8z�$C������#~͓�\��

O�~���<E/]	DY��P�<���d8i�H�|E���m��-A6唦Ӻz�^w��y0.��@�~��5h�`�@���VՍ��/�/6R博�����y׋x��#�3 ��͌���Vz�����#�}���4;�!c�R�TD)�.����	��-aL�g�^= "�y[��I	�Ҝy(+�z����d�Cl{Ֆ�F(�/_�7;r4M���$$��3h���1��L<u˧(t�oe@��a���ٝ��MZ�F��A�
ݗ�{�R�W�X}Ƙg�j��R�u��k�1M�A�ޯ�0_?Øz!1c�V�"���v)��?z0������oЀ?l00���'R�mҔ5H[���*`�~��>lv4G�1q�7L�叙(v����3_�o���u|��?~t,ț}C_, �sG핻��g\,ʎ��s�ؗ�8��p�r��&o��2/�u��'���o�q�T:zY��f�_��c���kN�V(��ijT�5��'�"4 Q��*���\�l�B�y6�^��#EV�H¯j�����g�Y՞���U��;����\��<�����]'q����yĩ����݌gsq�(�`�J���qM�MI,�h�N�ؗnD�Y�ln^��(�i�����PBXX݃\���b9����I��ӫ|$׶K&�3�\ba����#e*��7Vk*-5m2 +��}����fc>����U*f`6Y�"����)��6�Z
툅ו��/T0�0��>G:	z7h08%�Զ�)?�r���{�S	j��LM� 4?HW���`_h�s��I@��Qs���i1sk�Y�Y&\��}���2 ��(�pRDl�܋�d��r@6E�)���7!d����r�S#x<N��.ܽJ����0٨���j�-8]mt�(�Th�Nbn������~���}vP��-����%�Y�%]�� ��tg#�ܥ�-���Q	.բi��>߫���Z�h�d� vW�y"nrʱ��g��x�ku���X��a��%��Ӄ���%�ЁXTV ƇP�U�Z���3��h��얃�����f5��	_�E�V�t2�P{�^�v)��X�?ȷ=�r
뫷[,@ Y�; �T���޴Gդ%��Ѐ�;qУ Z�+ܓ}4J6vP.;9LAS#.S%��[����ljA�j�y��q]D�)�k]U�������79����|`���J:��}n�r��.ט��[L��CĆc�Fu�;�+f���"��aX�^�� �+��̩ʻ�'�� �g�8�4f�y˶�t�?�c�|�.i��(r�
��d6Y�܂�]��S)!���[d��M����p�ʖN=K7�Y
�8W+�n��%yLz��:�ϝ�����I�(��Z�$= ��k����m�q����X�1��r��ͨ����,���q�?��ȓǜ	Ks�|� Y����8��\Ir���U��J�3$�YЬ��$����('^����o�(�K�I]����x9��-��-&�e�J��[�������J�))���Z�0�+P�}��.��f@-���Gg��"�^HdVk��Y�|X�f��$k� �i;�Mk��OGj �9��ǋ Ӌ�%|i�\�UW$�?Yt����aZ�>�4p̕x�f�asҜ+��|t|)M�[B�q���o�|�Sļ��T/2�j�\}*���`RO/J�f%1���͛@��;�8����*����Ý=��wg�u�s1����f��Aɢ�n���.�IO����@����e�i3�e�ZX�����,,����%�cҦ�<��Hhn�In�d9�6`�z#�؂%�'È�-�F�7��ʫ/:��@��q�)�8/Ib�-(��:�J��_�o����K�#�!�uJ/��A`��vvIj��S���%�+Uc~Evj��d��c��ꌵ��>�t��2�����`����<Q0����`j�{|l�����zba]�E��!�:=�νSdKy�o�/:,�Ald 9�돦ٸnG��;k�� ��l���P���t��$����y!r�KƐb�yi�5���ю"��	a0�p8�u�ԡ���p���T�0��#�'��
��<K1=9��/<MJ��/\��^ �����OYn��o�����"v���[����Y���ef�\�u�}�l�A12�i�.-�t�g#B,ފ�pOdn%�ؓ�"u?������k��a�1���B�*�+���ð���
au�Y��|��w�5Tu��T]f�}�Jº�- ��N��L���/Tz�њk�^���O�{�%e���p�S)BH;% �<ۭ`5�B�S ����Q������mx�^ǉ�����E�3���F5�*�C}r����bC"�Zs'lȁq�LC/['��?+�u�0���Xn�:?�u���զ�Y�S\N'���e�2�Yv���F��n><^}���O3�Z��]��	���+'}�G�5��{p3>�Z�&{g�Z���|���mJ��^/�p;5!�
%�}�g�`�"�7��HgkÃ�D��Zk=��Zh}��OO�˫NL|T�뿙���������8y��+��.����k����u��AK�ˮw���B�3�t�y&�����8n����ϛ�U�&�����ǢN:��%xN	�n�%Í �1VӬ\�� Q_9������U�O�m_NGӏ�[�vB��mJ�^��@Ң�K�X�1����!��O�B�S���"P4��Z�O�Vf��R��{���*����ߢф�
�==���F��&j��;7X���#3�S���UK����gS��%yf��$CѦ�7����������\ � �W����ޙ�������A���c��T��z���_�vK��]ݐ���:��n����Y�(���k����sJ�rͲ�����t��j*MJ\\��[����׸�^�.|��
��6xic�����p�#kp����][�V�H|�^��]qau��R�-��nUWO�P5o�#o�zm�.P���Y�Թgz�Ɏ�j�_a�Z1��׽����u@v�@��������H��ck��W.~;K+Y�/�l��3]jg�=�S$2�D�:��+�I'[����H��S1@�ѱ�k#�y���7A� �@kbN�6��:���ϫI�F(��{K�q�ڵ��)vI�6>�<�%�?�'=�cz��܌�p 1�<c����l�K����L�Abꑁc�'[w
��5q�D�)�E(U��像�[3p��|b&�~'�r�GQ�g�{O_4��ċ��f��P䰿IS��W��ȱ{M�Cʟ~D3K�0�)ּ{ȍ��,:�'���g�Y�rzR��ԇ�6┍8�A���z���:����mJ�&����Zʺ�B~۪���=L:<*I�z "0�"g���oO�~-ɥfw�csQ3�DhOʰ>��KGX�`��P���ZY��m>re�lÏgD4�7,����0oee�Z޹Mw�2�q�,N#4���6�3+�����O;���1(���)��~v�C�UL�Cj��gN>�ݾ��}w��)y^���QD��L��s����D�z��	�������rS|m�flC��_9�B]�+��Y���&���+r��&8��ϫ�}q�q��Ag��a��3�⛱Z(S�����r��p�9e�|M`�@;`�?����B�Dg�w.�A2�d�,'�J	�e�D*��wbT*45��z�`�C�{ WSRЉ1k�b�#��zN֨j�g�R�ȮR� X��=5�ed�;� �n�?:����=x+�AU�h���ˤ?���a6��7�*���!o�lv0�ۧ
0�)V{�xn����%���?�.xbtӛ� 
%.}sAN��k�!������p^^���Į��EYC���j���R�7Z<?��:���QK#3��-c���}Ѐ�rM%6ȑk�� 7M�����0HR�`(�[�"�#���-�Ε%5������YU�K<��n���,ֳ�|zp�\X�����6��jOj��R_�/$X� ����eA�D'//<���$��l�#��ݳ����C��A�C#D�������?�qD[�A�����xK��k��1�O�է�̲��Ջ�}އQ�e.Q:�HJ�Lx�|`������oT%{��C˴>����%���6�Ꞇ<eY/μK@����o�&ce������X��i�,	m��k��}^�h1s�K�n�>��М�I�]k>_�$���y��&Zp�;��#�v�o�+�����p��0�`�=B����������qH]RK]��_>O@]��Y�֦M�ȱEN�r<qi�:��Z i Q6��lX�%`;np(j�3�M�����/ii% ����il�Z��b9��8�f=�4hD�����<���:����Ma���!a��W��(�л��gV&NEs�ΏZg���Ż�|�˃�шj<�:�U��1I�aH�퟿,���Ԏ���"��N��w�?���\�h�y`��Lf#��m�*�Q�^��ngq8K4/��������t���;���
��X>Q��h��JZ@&�y@ܯ������ӆ@�H\\���%'6���5'������)�D$1����!�v����=�IH�D�h���҃����B��q�B;rQR�H��=c��EƤDdo�Hz�.Q����\�A��N�[{�¯i�۞�;��(���E��f}��vL�^� �0$���!�z$ �O!�Օʫ�T�,
�Y
C^��wۀ���O� ^�e�e��b��/���m���l�l��μQ�L�e��Ņ�ZS�ev��Zq=���nR���x���ݭ}�,����� '�R���CUPb�ã�X��5�ئ7���]�ρ��m#=0s���`�������������s) �o�K 2��}P���� &i:�����j�p��(�媆m��m�^���̃�O�b(OB!�3�qV�] ��.*�� :����G|n	����h�I{ɻkn(��5�mr��i�v�����W`��,��cR�>*�k�'G�ڀ{��w1�r�kʟB3�s=��*w����� d���������
�t�y;mh����d]��ٸ��������-Q�M�Q1WH	�A�x����;�#E,�eDD��5��z��rVX�������B��ܛ'�'����w��V���}*�:io#֕���Z�A&���c�LV������}������.;�/С��K�}�Tr�8�.��7��M�L��(����'�vC|��#}T%�J��9a��H�%��{忥Z�Ԉ�Ă���c��ּ�[����	�`�Õ��rb`�^�4m5���&:�^���������7?�76�%G�[�m���i\h����X/0�E�Ը��D���y̩�ܻ�J�3:�2#�> ��Y���Z���j;DW����7�q��-��N�'c]x 8
��a:X !�(K�{̀,U�K9|ZI�$��O���8)��"��0�o��po~���c>$���E�H�����-p��^w���~{A�#N����ö���󢉭&&q/�����<�Q��u����C6���*HM�:��T��]Zx�<�h>���1F��`)��T�ڋ�Y�o�^|�u�I��<��ܰ�D^d�@>����c!�ί����r���Y:��cʒ��{�˔�=D��X�������T�[}�R=�" ^���bV�Y��~Xm����RD�0G��O���ަ�9�� �i��ვ�@׉S�n<���N������҄���/�U�ИD�NiȌ�}d�Ɋ_|,��1UL��@tF;'.��_��涴��8(Vz֭׊8u�<ꨅ�댙�Xq<n��Z�[0�XX؜�c��<8��V�c���w�*�R�@���2���~" _�
l8 ���_�%h�c �Hu��K����LL��
x��L��9�>?G]�xϒ��^X�X�B��W[<yF��	��*���I�����pߡW��Q��i�@���#�h��3��~�8�����P�jP���1ſg���Ʀ�򫝾%V�G���$�-��sӬOM7�p�q�����jL��>��AY
��?��z��"H����(on��#�|'���c	3��bL|�4ڬ>?�5S�eQ4��UTT�A��~��l��w]�z��'��mʈ]#��!~p�L�a�,��+�س��kޒ����V&�ꟀGiL�*�{拈�a�?���F�l�c�2��敟J����[��>:<�iR�&�P��e����4���99����&�0��}����������t�º�����T�Uʆ�MK�${u�Ø��@`�1�{J��U�&Z��٧�-�V�.ϳ��~���A����LNJ���M�M�X�1W�V�x�����k�Ap�có"u~��u��@7�M�,������j� }������s���=�Ԣ�28�#f� ��������J�9x�@�ğ��P�[���\�3i��hqr�2��wx���l~l�*KV�{���c/��,��F_�4�\�ތ.0�,��U����8%��I6�^��U��>�|�G��r����S�l�N�x���Fh��|�1p�*��X^�s�Q񊕈�=����	����\b!c[�����{���XU��2��v[�65�Y,����z|M�у��������`��p]���p�=�\!v�7��<"�C��}�<��ܐ�v�X�:���s��;���4�33�z�Չ�_�B�����=8<�1�}����6@���Y��x� �D-K��3����ދ���˵��Q����"`������ƣ�!��LK�C���{"O�m�҇���j��	x]�~wI�F���O�|�wן]�|!����+v����$ro��5��/���]
yCr{`���Y�I��9�˳��W^����0���|��2�o9�	�����D�B���T���7��iK_�t#�Kt��1{n�-E�O�Au9h���,W7/y��'�/=�����;�֋fB��u�,Ά�v�8��0Jy�T��ޅx|������'�q���r�IM����������*��t����}C	��I�H��[�~?���3њ��Q�Y�'�<��� �v�:go��W+��V�¸�<[JyZϥ���_Y�H�m�|fq9�b�0]�9Cȗ@�rUk��wi��U��SPý�����'�蛥=�;�B�		��x(��}	)�W���u��]�F��Y�k4���V|fu�}|5�ה�y3�sk�B������ ����0>���Ծ�v"a�󷫼��.-����f�]�u�C�����?�tS�
_����[�Y/G&�Yq����cPa�TA2�Ǫ�����ڕ��?�|���jT���.p�0弛5�P���q�9�[o�N̟��(Έ����~����=��3^���ꭙ�.�АKb"�T���a��w�����Ņ%;�\�LYB��"L�i��L潧Z�o�2o��8��|�*�ǁ�����n{d��&����}VV"����*�"j���+�����>�$XZV��s�?�96>��ߗ�2Um��]�:�,�%����������z�����c�/"*����+�:��(�� ���w柽�����y�tu��%��������v�����
�X���tp�[�'����7������n��:�PO���}+������x����Ľ�2��>�ۖ�ou!c�v�����{�!|�������M6�q�������Tj�Ԥg�Gm�������j�އ������CBZB��������K����n�z������l�>g�Z�z�}�g7Hg.��ұi�ӐHd���م}���=c�ՋE~�),ȫ]�-�W�u�NN��u��"8�h
��y}@���G�������X����IXO��JSF \�8�o��Jr,���O����0��U(�@��y��^s�T.�s�n��/S1�Svھ,gsqÛ�y{6��� ;�r���������c������X3�9��s��'�p�1p����36:��9:�F~n�jd���*�qWo&��nWp��]��S�+3��L��	�=|��]�>�-��M��]o�~Y�U�\2��)G����"��`���d��=�`oc����+Wc��O`|�<o��U'�!�� ��c}a��\�(��,3�g+h=���ɨ�L�I�w���(�k2�A��(b�FEj"�&T݌����c���F�ᱣ�cC��+K��4#�� b0nK#65���Ǝ����z���Ȟ�0����o^5獽C#,�¶�bP?	�j�R6����Ց�s�ҟ��4ᒐ�D��CJ*Xo�k����%�<$��Ƹ��+��(O�s�j6$�U�F>��.A�\s{�7%��yy�(�)l�=�B�=���=���y{�e-AxrG0�Q�����k�*��a^�]��f{��砗�ܪ~H_j�l����lg%7��oʠN�����]��~�zywhs�*F7�:��wh�����d� �ϥp���Dk�5w�I���N��N��N`�\�n/�,�-V�P��6�42���&���o;�	�GY��t;�y8#K�8�	�a���.��&ێ�_��<�ir�׊]��;��\!3��z�l���ptG��)rI��֢A
�
~g��VBn�B�F:�L?�/93�$;�����dN���@ܿ'G�5��7c�=Mln��g�Gw��Ǽ�����M^����S���ɴ$�+i<.x�C��u{��:p6� BC]��LBFBY���pa����y{ȅԿM�]5����[Ն�M�������4�#g���X�U�fg-ߞjܞ�8[/�A��D�樉�$l�̐ۈ�m���r�~�����������6�nd�/u�z��߫Ȍ��6?�
A�['4��D'���e\�l�:`��܂�����Dl����|~p������D��[�l퀻rff]�ן
l-���s�`*�����uM���2��I'��$R	C`��d������֣7�_*`@�6GQ�e�!i4'_6��(d�֓96��;H���S��N.] $�	2'�@��4�18O�W�n��T�	0}XNB0_��@��]0�Id�n�`-�o0�`Q���+��J��U<<<��)H�Ŕ�uY[��fw�}��������R�Ep�D��).��}���,+)=D ��v>�b
m,�p�'kp&h�-�4�0G����S�hmW����>��]U�wb�eb�����K�Vפ���{��Z��ͼC^�H��"i�}�$�;t[Zc�u���<˨���ͣ�Tkzkw���'�{!D�-�ďS�ꪂ9��D{t����o�9�̊IΤ���[Xj��Nv�d����x�۷�]�ɷ�	L��K��GX߶�¢��r�M
��[@tM�,"�-��a۵?�!�R��Hd�yو�:WO��8[��0�/S���ъ�,�dE��T�*���YBrYllB�h�./o���Kt���ۣ�-���T9x���'~��i��:e�K,� `�0��0�tȞ7=��m�vo~����O��,쁙QUkc&�S��E��������=YHR�
���g�n�lgoP�w�[�@�ɲ�B�������Ê�%�(��6��=�k��jg�V�l��K����JY�H�{�pp���C���2�"m��a�?w>i�xq��D� �u�'UB���ձ�L)�|�W�Qgs+��+Ԛ�L7M�ə�yD��,��/-�fy��O�|��d5#[3h�D:��U������	��+m�@,(�ѫ�?q�O��y���E�30/ �������BWS�Kq�#�07fhfUQ[Aǟ빧��7Z=��Y~U����IԷgaA�x��w�9=���-��w���FD ·2��4��so����)B5�R����	�'�cӉk����3�<p-��|k�=_x#�Վ��7��Tٳ����j����o�ShT���@_$B���|�06&����Y���#���>	�t���0���n��>���O�6�Wa�0�-T<
�(��}gg�ӵ�C������H�%|��j�ɿW�P{���N��o�ה�<�;��u�}_�j�]]���{�:��l��ν���F�׮�ec>���mӢ�O"gy5K>�}�`�|L��	��0�s^q����^^K��LY����Zyj�]|�O�^�w��v1q��'k���y�Qo�v�s�n+K��МI� �DQugd�F�����"��oBh�9�M���UR;�j2.kԷ8E�;p#ր]�.T�j0��E ���}Y��'[�Q��P���A?�G%P���c!�{`�nwP��1�&���{t׈����)��E�/O^֏`�?&�>7M�ea�y���J?6\��[�e�2�,�H ��5�;]�����/_6�,��ڮ)J}���*'6��س���N>�����0%Lz4ʙW�O�ȵ�>��v��d�@?B"����4�|�uӏk���6�b�hw�$[@�y�}�g7M}v�,V�����tQNd��?�!�ct5�w'��ZX4�4On�45��ka���@�Z�#γü�á�~���Ey4҅a,Zn�xQ�6.WA��?��L�
�d�A$Ғhv�� �uO�3y��9���L����_��Ĳ��F����=��ҧg&-�03����K�ӎ��| +Jq)ۨ��
X�u����Ϟu�hV]���ă������1\�Wl��@�!v�)m���B�J) "vMu#Xq?����l�fFZT�;����)B�"�����)}$i!�!Ao �����7�l�R;�k6[ݠy�Y�8��VEV^z��i�����7�U�@L�ټ�� W��.p�:���p���J��K����]|�P
~��N;(x `�1�ۊ������6b�;;��S�Mr���N�p}b�%N	�M��	��	�&��b���78��n0��=�;i��"u.�����e� '�[lR�D�R�a�F�zr��9p�����ד��U?K����>��v�:,���B���{b@��m��,�?Z�\Sߑ52C���� �ʼAc�8�F8i{|�X�$�U��d�*Rx�\�cY�z˅�ADozcǼ~;{"j��Ʌ\�8s�����7�K_3�m�q�b ��syXOl��
��!t����`�����#ܚ�/:�~s�^�����6�������wM}�W���+�L�_ฟ�DK��I�ڝ�2�ǃ�nb�2��P�����嘆'�_8�~���*�G͆�FYȸr��Z���p׳ċ����٭��C�8�?�2D>ڷ��]i��V7�������U`*�Ɖ�b=�->X<c�ւ�ر����p%���ʷ�kPW��\���1v$)���wj���G�����yu��ـ\BЕS�(UM����b�Xzz�7Ooiؽ��!$_�n��@.�"�X�\x8|P�:^$H�Z�����w��� �;���
���\���R%CZ�`X��-�~��{eu1�F}�H/1��z&%G���uh�����b,ZF%�`�Ob<E�/�e=�J�����������Nͫ�;߂��ƞ��+�߃sUԽ��K��1e�v�����"A��D��L	���(�j*P�T���m��d��P�}r�YFY�#D��~\��)I�tFU��slF#�`��m�h�Hx�^�(ke_�"��g��o�WVĽ^.��0�"9��7� �-�H�Y���$�*â���{.(�M6��gv��2t_�3?'����DG@��ڸ�j���Ȕ�m���S�y�Y�O�շ1�D�ٸ�A\m�>�K=�� �/s�r�����/��j$ow��:���0��-
�,6�&I�+ �-ߦ��уԮ�? m
~�F'��� ��i�Di���Ĭk~�{�7��O��/� _��-��;��z)�fu�	����H;�9,��	�{����Y��.�����! +&�f#ؕ�����9�Z~�����2Hfd��_��L瞂�
k߀��(-�5��B����]ٗ^������$��n.���W����H�<�������?3/k?`	h�L�����Pey]�UN���N� ��vGO�c�p{��@^\gȻ���&�oU9ʮH>NIj���`"����j��΄��	kňj��ͲǼ�S��$� ��q���*T��oŶ�ZT�@e����S�蔄�cPh����vnET���J����9���VX�M��[�J/:�ՠ�J�w���!=���#*Z����ץ�.];Olf�7�!�l-�pC� Ġ\��C$���m��g�c���c�7K'ֺ��R=F)�PN����:}���O�,a�TvW�UN~�%�F�����{�p��:�My$�FI)f��p��w�-$!����ɧ}��̊�à���(���E�AF���N�ICc�3|��"-;4fC�G�a���s$�㺳�s3�|ͯxݶ�u[�A��܏���sւ��z�'��c�Ľ�]�d"�m�.�IRS��]����C���������^�.Wն�2)7�yp�L_c��A��_��ԇ���G��PB�?��پ�#��s�9�^���[͇U�6~�m�R'B	hJ|~0I��
{� 5�k�h���"��C�#拧'
>i~L�
��z�>ilM�?��+���I���h?�!���7S����R�6�'nK>4�IF/I�gݹfl%`:�f�T<�W��.�q�::r��"ϛ����PU~���P�W����9��3Ő���f7\U}��h&�x�S����N����v
�y��;�g^۠�,yl��`���ʸv�dK�s;�h���������K�Z�#_�=���I��|Ƅ�N�1�|uC�L�5��ҀH�@5"F�H��DZ�{���9��h��,V,�}]E�y:E��������7�y�'�WB������OZ2���˲3R��B�/o��W��|jǝ6�1��<Y5��.����m���P5Xt�����p/�{�d��TWs~[c3�I�"�lUM�����Y�B�99� �'�[������V:�q�`�\���08�A��Lr1 ���R��{���ueTٮd��a��w�Q�{�<�a�0�zq6�R���ն�=��֊��PM+,��&QE)A��L���][l7g^�4�O�qC�ダ���*�ߥ�������n�V��A���Ő��ެ/�5D|a�_����L��8�m��$�x�d;�yh�]W�t��r�<A;��ߺ�ʧ"M����p��&W�݊����_
 ���G����a2�f(��-�2�z��t�f�.�_���r�4p��u4�/$Fo`z�S�U@��B���U�&ig�y4 P�n�_�u�Qc�W=n/9�h;�6��Ah��X1Ga��M��]�����^�)��kWH�Rl23YI�]��_�)�q�A�-�3��n4W�	O����z'}ї���FV@�]�F��1�Ms+ �<�����y���E.�&s�{�b4���p����x�����n��ǰ��A���5��oY�@�O�/-[vP�tҧZEt~�-F�3�Yz���@����_݊֩���Nt8rK���s-92)j��.�������%���<4����j)7B�k�\w�o�y)EQ�S��o/b�4����fYT��k��E:�IY58\�����|Jn����`M�G�������2�(Mb�ț�G|���F0�ϳX)u��_���
��;�;:�oN��|N�R�6K����w�ܤ���=V ��s"#S���hm?�~�B�c���s-�M
�0X�A	Y�F�#�6�I�T^s~��N���$�}� ��e�Q�%
�߈���}
���0&]l��_��o�ѯ��1�* �1b�X��u%ō���90���?Rwf#)��S%ʔFbڡ'�Fm~�==fb�0��PMᯡ�'㷹��H��F�IE�탓|�fw�[�>X�[ۼK&��`�
Y������۵y���
SMq��v��eo]��=qPw�{��Ğ<>.��/
Rf�v��vms�����*�%ƥF|el0\_�X+��-��Z����:꥝�˸�E���f˾@�7�%ˬ������h
F�U�D��\��^����l�`Q�l���%u���lAۦ��F����}�>��~�;KL8������ oto�*}��-���@��A�vm��m���}玏���w���n�K��)	x/Pëg�u�q������hB�����b��w��*y�\�ٟ��)(3!չfSƄ�u:�j"�� h�?��W(x�|uz���w����C'�)B�``oݺWc��X���߳��<���������P�
���=��/_~���F�]�[�CiV[j/��u\�{��3X�bd��.cP�R3bM��V��K�6�l&�>W.�a���wj�1�ֲ�����LP���f�vt��{(���aHr(_��Z,�9'E؝j̀��і~k��t�+�89��*Z֙~� ��͌@��Xo0��E��X_�������D'ڼ9��c�
C���ˮ��M�ޫr� �C'y�M�1����i������f�	�����7&0��{p3�L�)5a�wu�g����3H	�!��?gҘ(�q`�R�ɇ�5�27|���)Z��P�bp�&4'�V����C�x�/�5��lX��gS�`W���Lz��
6��bQ �4�z�T�����@,��TLg����[�z�PD��%D�%f����ڵ瘀n0\+g��<c�l�������%�7�~N��A(351d���.���)Ӂl��DaA�/����Oy�2��1ƾ,i��2*�s�W.KW;%3x���0ơҽ���A�%�O���TdG6Xs��X�H�,,���ڂh���v+�!��l��e&�%X��~�_��� ������>�5���om����n�%4Ja�P���R##d�6�jG�"*�$��q��?�~F�a�=��wB��X����GK�(������j{��e+�:��xV$��i��R_���w�]2 ;�d����;d���\���[�]�u#.�m����>��ʇ�I�PQ���5{�[T���=i^�KٕP��W*@c�:���mU]6�}�ۮc�i!�W!��lB��C�3=������ǒ��O%�����m�vL�ؑlWG����7S��^����3����)|�Yh9�c��$���[�&P-�u;ݺ�7�R.��E9�@N�� ��L̃3ϧKU�:�����3���N�a5�'�"(�e����OL�����H:>Ó~��[[��f�Uٷ��7��H�Ѐ�G�<���▙�Q6u����p��2�'u8��1�;�����f��e;��p٧$7�hv(ӈ�X��^1��?��:-,��"*U���Y�u�ܐ���fm�Et���}@�T�U	��|*~Y�A$,s����lGf��t�j�u�~��\I���Kt��-En�:�'��\�����c����m��J��ã���wM�u>�]�2(J���䜷��4)�u?���EZW3�]���W������_t���eQT����������}���c��ټ�uؾ×w?��#��j��;<\��({����l|]�����/��a�*w�^�ႇW`�H{�1�4_��0 b	�?V���I��#O�u���}��F7��^ui�����
8�T������hIy��Ke�mQt�_/P1���Q�;���j���K����}�n��X cCㄮ;�(��)D��cSr���%r�)�	S��S*Q�mMd<�����׹q8���q�r�6xx�]��z�A�����7���8
Z�������[k(��_��W�k~b�f��+�,>�2�hWU��_h������E'u���Ht��u�2����7n����y�Hf����Hbݶ_#�F0�o~�}��i'���~`Ct@[�Y<R}���o��u�����2��	o��䩔���+�qjޮ���X��๶9CjLk�3v$��L�s���fWYy��<M�oT��n�I�6V���m�nş�	qMvS(��g{.P�/��Q���?��#�%zN�K�����!y=K��q>��1�<���}:}QR��X����ѷ�����I`b�_�"h�"MW�JX�8#fd&�o[�M'L�bR>��EQr��w�B�,��r3ʁ��ugv��^�)��:�b|ڗ�Z��'�@�1t#;aF���ê`^��P�D�����8�l�2�]HqWa�ňQ��h*�� Wzm<��<yd�
���S9XKɕ^P � ������C�Q�����`4[0 e�o�hj�n9R������v�Q�"���8��}�auT=;wd�_@GM~��W�3���^����<�}G�%�מ��YO;V)Nj� �����AqPڥ��^�%��9�3.)3`MH�������A�r_(Ťy��-c����������K��bN��� ��� �Ή�XG����g�垉��=IJ�:�D��r�� #���1����<<�������2 B��_D�9y��+x��CG�9���X���͝ɲ�<���_���ۻ�C>sb�P�9�bp��j�'f��Q����Ic^�z�����{0��Χ8�fU��҄7ߧُ^.�~p��\=�~�3�O)t|$��FMDfV�!yn�M_��P��C�'���w�x���u�k����(ll:�@^o�z���O��6Ul���)�g��W׺d��h@\�"�@��@d�{F�\�~�h�z�`��(8����@n�~�Q���M����G�q�\�JBr���C���~*�?+�� �uW��g~p�&�sh��_Z,�`������K�W�h��C�՜�|��;��ěg܁+��jQEU��r�Y������^j�<>�2���݈��~h
I�V&� "SRE�g�%��Gm���a���Q~�0���+�!�����K� y艡�$�YG3�P�{��>tdGSC�p�;)7�;iGE������5{50�@��7��hG�_����{���!������1W��w���>�|н�&RWJd	eJM���d�?��K T9'Ņ���-�O�*x� <�-ҽ�+"��s�A.q{��r�{M�-P�	�O�y0�I�u���i�=IL�}v򢎲���	���Ɨ/�P�!�@!�?[�M㹙l#}>�`U�~�$�Lqw�G�IS��] �Spg)���A�c۴��p�@$xB�����ht1U��:@�����#�*����g��y���k�DB�+�l�kx
C�T>cqܰ�Sd��:�eB�v�i���Ƙ���O�ȟM����3��ڷ�!���J�q-&[�[��Г9��TE���i��* ���D�{T���ն#�ҕ[�@<���n�*�8��s�m�����B�2�pD�S��C�lf��a9�,�P}���C�0(E��:��ˌ���C���5��Fe����&�_z�R�e#�%�I�ք*�v�+$�S�7e��ۘgs�[lvsD�i\��6���{OO���5�\!@�Q�T-��<�7-*��n�<<���Ud�g�����)̀�V�,�P��|{>�I�f)�(��ϟK;������B��<}�1<�9���D<|�0�ؔ�'�&�1��0^(��?��.Q3��˩ӂx��=zh�2���4?&��aL��P�?�PQ��o��`�l�L���D�A �[�=D ,K�,��Ds���>@�ޣ�`R�����8Ƚ���t�=;����\�R 	�"�F���EA����<�zLY��G!#a\��
O���j�=�Ӻ~���k��~�ШΘ[a���z�OU-�jY�;${y�ѥ��1--��'_��X2)>9),�k�%�f��毷����]X�𱤫\��y�x!z��l��
��b&�y�e���L8�l�Z4f���3�D�M� �E�҉��Y(�\"ͳOz��#��ۄxԻ�����Ӵ��C���,M���<UX5�%O�ڈ�lo��UU��%
T���7��������_�y�yPZ��$����o&�WvN�%�Q/�`��O
�����U����x�S}0�so�&8 n�R؛G��mz�oOSyND�7�|�a�4ko��`�����)R�ǰIˑH3=�p����R�����ת�xmm��� -Y����� P��>`�0q��0ڒ��xo;�V���զ;�i'Pg����ÈG���[1Fw��b������%���/��!O�q�*�o���u�
��+�$�F��tH�گ 1��X������?_T�'��`eR(�ebSq�g�Z�nF�y%邾�����C&x���kU�����ܣHM���9B���i��*.�*K��s�dЖ�\q�ڍL��W�����xa�w����L�����̯��R����N��������5��s�I�X!t��fU��2@�Cm��sN�џ��X��x�*KO�3� ��Vi9N��� X��BOa!>j|c"�}&��if����5b�C6��j�ɑ���=%q1#6�˲�Ȉ�S2M5��H��8���	��?�AD���u���'�,t�&��`Y����}�:���R �W������q�<�eeG���R3�����l:���$��$ٟJ0`'�����	&�0=�ⳋ4{�@�d����&�u���.�-�/Gz��K#.�rh��",��'��Roa��?�0`+x�@�w��&��r����;D�h7�Ę�����{�I�����k��Vb����%�ט[M��7$�k7\�����A�	h ��D��F��.b�#�gu@��Gx�<PC{>uxK\�-ፎ�*�k���;އ���]+0��^��8��,�`;X�qi\��/�Q�̶
aRa�X����㍆47�Ym*��H�KW,O�zY��4�˜�H��^g���A��<��)�����J*�Vs�}:t�т὘��e���L1I�D�1y>ܤGK�V���ϩ�2�OCP��2��y��h4�1��J	qīCf��D�Fv���`�a��	pX�} �U�q!�����LZB"�$�f��?��<�8k-9���S��9GҪ�Ԝ7̠��C��p��.���6Г������=�>�p��RQ��7�g�e�:?���|"w2��h&m<3`z�q���:�B��(��c|�w�Qu~R���F�7�L�[6�C�`���<~�0f�W�#h�iy��%<2�9��L-6�u��F�pa�h����M�] ֪������i��T� �z�� ���B�coV��Z���[U�k\ub��/�HrA�ӡ){QSt��ZfP<����T��1�{�����`�/5K�<�G��"�]����,��s�c8�'�\N�pRu-�x�6�����Cc�O(�e��/ŏ8��ZD��V_ߑUD�2��E���".���$N�A�t�j�)Y �_���՝/�&�+����S	٢����g�TE`Hv's�w�c��@���K.� �M�9�Z�T	�(��g�Re������!����6
�?+'g\�d�G�par�y��T�Uz���ɚ\�T��l�Hh�h�}0�쥝��ěol��+�v}�-��rz��6={顗ƈ�+���R���!����+��}u"+�Z4�<+SV���ό��7��eI��߮hg5{ϞJ���	ZҰ�跪Ȥ�� �ݡ7����;�-��?+jɌ;�������	'\8�Y�����5%��7o�.t�~2Mp�a��mB������nd
�F����c		\|]�y�jn��&}(�6�~���O�9�H ,����5V	b/q����$��9Č'���(9�E-�;3�+n¢J4��2�q[���&�#�YˌS�/_*��Y�aø�s�����i�[rF5�[[9L����@<�y��VZ6Z(P�M|)��L��*g7�2�2�WD��̐���8����Y���#����+��M.|��+�Ay���;����X�faE�o'^=�S��(�$�Z����B���>Ξ9��v����Ih����f�w�rS�3��[�2��` UUǢ>��GB\�m�zx����L�7l@f9��"M��_=�
hv�1Lr[��6  xt���7C��^݈�\b� E�Aj�4��ʨsy����.�S�z�8��oZ��Q����������#O����a}��~�o!����׺5$��Gb�K�����hk!���]�������� I���:��H�W�B��K^����>�eO����?�DKI��y�?I�m��x��� g�@'}I�	l����闁�H{�9�[^�<��V�5�c�C�T�����5/�Xi�3c�WU>�~��u�����[�����IE��I73��ZS�G�w/�+�i�y��u�p�"�E�N56�2��#�}�4 ��-�J��Ɵ~	{;��^>��X�?@��!_���|��@��B4�w�-�'�cm���B���+��HI��wD5:�.��
���7I�!Ϊ!N�Xԫ3�t��Xf�͖}�d��Xz��KHX��|Oˬ�� ��D	AHz������t?θ�ߣ�>h�\��A��<a'C(<A:ݏ����'	��	aj=���Q�N�~y�|`��'�-ޢ	��5�^���6�@���&U�ϕ]��JG�O<ѶwV��L�$8�����Q�ڂ������`g� '}	����̃krI}yH���i�Q�C�g\��27؏;ռ,�{oY �P/�������$���Q��1O�M*�*fi��7I_���Š�1(� g���-�!�;��ǻ7K���~��6�������|�c����m��B�� '
�~n��X��O����w��H��;�9 �'+�=>�y�+�'�d��0��`\�U�3���>v��#�õ�|��3f&��~��	�6��t����(����rT]Y����Q���O�ʁ1p�Z,�r8��t?ٸ��*A�D�G��/���S��!N��W��y����Z�����|̝���,i�x��W�a��h2��4=��߿?��ś���`0!����]�9;!�-���iC�J,M�MY�}����a�gk20C�������:���: �RvFH��:��eD�*�|��N�zV�dpP�I�,(�P�xKs�Sf%y�?I��-0=�"�!��4U�=u��w闥�ܣ��/���:;��	�Q�� ƫ!���U�V���e�Ɵ
��O󉦸��:��j�AS/(-���rJd�ui�c��>��Ԣ�IK�4;��	�;��j�zu�y���Nh���<�^��s�>] �������Yޞ6��V��D,{�$�"5
4@�~���p-�z(2�G�A�6�E^7re#
���)�ِ�6̹K1�O-�Hƫ94橇�����3{Z�@��޹@{⌵��]��.�2.��p>aҐ����aO��;��~�������̨6�~L��^2�*	�I��c DB#��Nb��^��(�j�\n�5Э�,�0n�S�qw����y5dǸ�/��GP'�W�&r��k��Լ�ϪE`/Aq�0 �_�'��c�Gu��:����'��%����r������8�u�br@���ׄ��@|/k��ƗRs�����)�;N!ۃ�x<��Q/_[�7��FB�@`�!W4������Mdm�Z���5���į��Җ��7�7Y(�99�(�= ҇���)3}�����y�vˑ��:��mN�觎����QT4��N;0�p�K�e�8-�m�Wf$�"�
�Z�K]E��/)Q������鰢I�_������P�W6��*%G�����Z0�������C��~����I��X��x3��tC���^�QCN�Eu^�_q���6�{��U"�2mxW-��og��p��750������ux	����O������Lwqeh�	��NT(����|���Y%��!��1&Ǫ����rp�t��m�=��/:&�\QXvg�AC�/��;����|��':�4�#�IT�i�J���w�0���f�N2>_��h1v�]�J¶�n�9M���{+	�[�#I/��c��X��a�4��$���c� [-�N�*������)B�Vf��Wn��aAg����֩O5. Eq��J.5��O����,'8�f��A)'ZX��U�	��
uƁX�F}�>�]��R�s��2w�7`�5�������/��>�ͣm4G7N	��$��x����w�`�e-��ܮ��<V2>��8]���f�vx���p��x��'ֶ�x�Ś�8���Q�9��w���i`>��iqH�/.���p8[�jVE1"�L����.�
U�(�O�B��u�����8��=�2][gb�����Xژ!?W�^jv~̰�;v�ŏ^�z9�''��-�sb2�[�;�VT��C�Ҙ���Bƚ��yq�MXU�u�����|(���ok�������y}b�Uv�׋�r�%�v�(_��eη�4�Ӷ��C��^4𕓬7\�D���r<r�,�p��Y<&��A�VS��V���]ay��wV�k۠��SI�?�l��3��	�5^��Z"����U^%��k4�/���q����q �}a}���%�ւ�߇�E�����ռ��c��v�S�M��|ׯ���9�`z�$2ѱs��|JJ�@0���K�H8�����|��#����x�OGó߮�G���4I���{��K�gX�?��~�1�_NmA��2�d�����c<�,-�x�7Qŀh/�}����u�A�y���)�K(���U0�V�#g�۪�ͧ�"�4�Gٯ`�����T��$+;��Z`S�Pw���		ko����Ys�<L��%X��ڗ� ����H�8ןA�
�/-���6�����oD@n�������7d�Lْ�ZJ��g�8� 6o%��ퟫ��fDq@2�KD�u�Q�]!0Fqz��x�Y �͓��f��I<|lw������_=��r���d��X�%�ق�r�Y�T�"<!�2���4�Q���������5�6�?�$�z�Ď\�ٮ, ����=������ ��T��u���5Ӥ���8`�fz���|�n���������7뀦��T�Ƥ��.�
��xsi���e���XB,�{R�t��5�o[���t�%h������I�cf��Fw���J��۲1P)�>�Y�X���Y�+� �.��m8��.��k$ߵ�����}�L�)�\��}{�����Qs�����J�(���I��׼��-��Пv�Ҫ��vPP8��Bv�`�Q��j^�!9P>B�6h�B )���%6gI��Ff8n����	�Ň�rii�����s���C�}�{��m\���K��+m��.�SB��L�ڵ�[��D����n��X6l���9��nO'����J�q1��\��F��CIy|~����)���4f��*衂�[��2��r�~u�|������;�ujy����Ǵ읕���/XDD����;U�+��_��n$�S���vv���T�����X"�O��鈬o�74�E_�V3����x66D�`���N�*��e�J���+1³7�dFe�O�K���Z��H��/�Ff��6��"�
j��\�*�bI �l>���o&����w��L�b��6�z>9�����00�#^�Kdґ��n_�:�ec�����ʲ��!�T���w��Q���]R��b����e?;�m�I(�������H��)�ikU�\�<)����t6x��l^T����0�u� 2B�G�_\�u�w	E�v�FD&�"�
Ƚ�H�V~�:�h<|�7���Bg�}S�L%fe��ܤ�L�p�_:�=#��J�x�&����ZL�ߌ'���B����W� E� 3*�ﭥz�M֛XQq� D
�7�r��0E�q����UJ����Z��<;OG!F��cVY��B&��f�n,N�B�ϣ��׳.��;����澸�7Y��v;�������O
M�L�^��)[e��1$����1�ra�G�i��*�])��Ns�2���e9:���C\�����ԅ=�+G2"w9r��F yUQ����p������?8�O�Hi؞�z*�_�b��&7���R~4�9O
(�_�� �L�!�6*�h�����h�g����?�ڶ J]�f����g�LO��v��{Si��@��OU����60DI�~H��\���I�u��^c�.�XM�L�$�qm��5w|�[m�6ak׸�R�}1����_Q{��������͌��2[y��-��J���&��f%[��b�N��7��R�N&I�.xH.E5� �����~�E�c�"*�ϩ����udcB�%B�U���Z�?�Z��5�Tj��4Ns8퉹��U�m(Qy�5,:��]��\lp���p�,gC0�amo�y��[ϰq�p��
/)g+􇙔��"�J֪%�gs�K��fKU�"���K�}�#�I������u�D]J��V�e���?�D�(�W9M�Q���Jq݄��vי	������\;��3>�Ə�
�w���U�G(��u���C����ׇ�V�r��(�e������0�3�B��AeU�|�g
E'��OL��_��F���=i\�ĝ$�[�hC�u�hM��KY�ڕui����J�Tie���V{�
�u)Bu%B�"�6~�U�:��r�|���}f��y�����m��Kk
�գ��B�~۾Գ!�fdk��4=��v"����9{�+��by�F}�l��x���C��.(��ܸ�
O�1ݚ������w�g�`�?+��Ƅ�����>�����bUb��!� ���QJ���[�q�Kb��[u��Vp#c�;z������+���W�����ͬ�S��_�±�"M�C��o������*0�sw� ���j�v�-����>yMg�n$��|⃸ti��S*i\��/���`��ڵ�=�����g�d1��]�˝��xU��&�MG��|�d�>�+}�ǃ���b�ya��̴5��%�˟�FR�n;E�#�v�3}��ݚJ��Lc5?��V�@�xP`����-<� �`WQ�x�S��xw�M��sA�FV��&�x;C �*�*�V׳9���p/\)��ƨ�)��#;���q�x��v��z�K�u�8�����I�u�׌����d$����z}�i��+{�ǁ��R{E~�F�5�@,�N4��i_�ǫ�о"�u|WR�dM�`�I���`$)�B�Ճ��t�\�^p�3y"+H�9τ��4�n�E���C������Upm�ѠQ��U����ifru$-���f�Y9o�g�,OKa��`����-��L[i�c���B�=�a����3�{6� ��p����+�r??,��=wh�z�c���L�Gf+u������A����zKP�C���A��Q��!��x��f�qX�5K�<���/o�0���85#�ԝ� �����S۞����8ɚ��u�-q��1h1Y����+$�c���V����^�d�E��Ñ�.�PI�!q�gԥ^����'�V'���#m*��NWC^��[��!��#F̙�;�w�$��mf@>�����y(���H�Q�U��*���Y�*�YԮ'L�t_q�yЯ^�,�Ɖ(��/�F���P��Q��3�m�䮹�o�}K

��*�uQ��2���+L��WN�A����0e���1�٬Z��"�cZ�n
J��g�R
�����F��B�����o�����\�XM��α�e�X;/��c��@���O8�ic��P���(�B��+;�ʗ�]7�T�u@*"oG��������s�\R^���̲-�8.��-L�GeT���R
�ˋ9Vs������Ŀ���:�d!�kJ�u��q�E0���.[�Y/��^/}��󮘾�R�ܓ��P�V�~u�?ö4��5A*���Ɍ�����<��Uhj�Y�;���*���)�c�X��1�U�����Z1g7�p��#�1��U:�C%�N��5�(�cȵ��񦰈?�ӭ�w�����������䵔.��p�h<��"(/u�(}��
G�g��T�[�I��H_��7�A��WlK���O��,*Vh_�Pih3}�7_�LM�t�hZĽo��)�-gI`��?O��W�Xf������^V���B����S��j�y,<5}�W ����'�Z��+�ψ@]KK��Ci�ۑZњM��/��*L�r�>���M S3�G����	����`d
��P�O�$��L� ���4�Ó�3�I@�.Α-S�2���i艶ͥ���F�T^Y�MtOL�+T#~�	�W�����!�P�;_�7��~���]��X���5p�"�>"��<�+����i �L_ظ�Bݬ2�v��ٳ�[�ޅ$�-��̬7���5X�~$�s�ʓ�C�����y���A�Fn�e��2����,JI6���.�
�t�Ø_�����0�5Zd��θ�����`����<�X�<�
PN�i�p_?�WK��~x��?�qO��7�P� �������oV��'��=�Ӯ��_����gDY��%�|��#��c� :sv�5���0�e7��F�%�|��kZ�)ʘ\�j}I;z��RvM� �eQi9�==�Ǌ�Zym�ˊ��g1gq�y@�3��c��t#�Ky� ��oٗ=0Mq�w�MY���ݩ��L9�"D�m�>3����[�~�8�,�M���^��Be=�	��'�~�8��F�D����}U��G�_�0>�(CJ�j�{�Ǯ��$��H�_)�V|����yo�,���ԩ�0fT��`J��w�	w�¹��u� ]:Q�뙏�ޛ�0�w��X�����|��k��	��%m�@��)�W��rnU�ӷ��¸��m��]���ev�8/��2��«ǰ����S�pK�
�q����f��>����%H!-G!�����/>��ok�M�xt�՝_�~K$j=(�PK   8��XF �.�m p /   images/9fb635c6-6568-4694-b870-d787cbbccb08.png��T\M�'��Cp���}p�$�;Cpww�5Hp� ������l��}���ݳ�o���=ӷﯫ������T��(�`������`��J~������n� ���I����j/�����������RM�ISQA�b�fh12es������D����M� F��v�4�MP���0��"H�^���R�����������1�	� �&������!�����Q�M��_|����� �q����@SQ q0𳱳�@� �?%.>~~ ���rp�r�@��܀���Ow&f$����ϝ0����� �������q0����A@�?VGw;'C7V;G�8H�:;X�;YB� �A���ih�����?l��������l �?@����l�չ�1�����������?X{�������?�����DQ����ЎNR.N�=�Q��������`l*��g��5��p05t�8�A 6�̔�?cpp�q�4,�L ��o����.a�?���
bg��Tc�����d�	�@��*BL,���OPnv����fL���`c3�����-m�M��v�4���Q@bq���.��b��( g��dhgl*')L����D ��m�e�����o����2d�7��g5����s�r���^b���������g{e�?�eh����/��'YK�?����=4��w���/+04�˺�i��5K&4W[�?k���]-L�����7�b��j�`*f�G���9��_r �w�����S�'��O�s� fj�'r9�	Q\�6x00��r�bjnG-��&�Z�)��j��7eIS��U��xn�FH���f~ZBmbbg�H^�����5wTpE�z���a�-	�f~�Uˊ�4i�s��h�?�+k�Q�,���e�veD_�yY@�,K�Q�1�9_S���cXt�";<<��q�!��8⸠����.?���%.:$:���zAn,nՆ�������Kv�@��_m�(����|0�%5�	g4����73V���\�����ߓ<��v6_��{�^w6d�>�?{�:�/�雲��-��Dޛo���/�8���;«����Sb�M�2�t�����;X���j�ulW����8�K<��q���+O��$��@ߣ����	�,C���=7V+�;�'�)�P,�������/��^o�k(���'��P��6�SJKKM��t� ��N�h�T�,(�(Q��%�[{��"��BT�Ů������_2J�?>�<�_� HFs��L�.�r%�5��=]<Z���V��[���:�+҃��/�)[�[��VO<j�_��.��Ʉc/�n����N��r����X=p:�&�@��K"o�U��N3�9�@%�%����0e/>G|r��ljZy�~{pp�y��R5C�����kN��#�\��g�Ϩ�1'��t���T���4�b6�J��;_4�L�Ǖ˄�d�N.X��������[$c���=2������~����vSb_r�+Ӡ�f�:�/��y�X��8���٫�A�����Qd�{h>K I��}�BZb~���/���3J�͎p�
A��S��X�_vt�5��7��ܟ���AY�ٴb��?��3����~�2h�t�S��ē��e�%�-�7:Cv�_R|W��Zy�܎���C"��j�K����c�E �y��b��"-ӷ��� 4d⟽eX����
L�"���خ�_u�]�F����������5����"�j����6�V˳��2�޳�����RT�c�u��T8j�Q(Sq9�Τ�i�����w�*�8q{����ٖ��`N�#��u ��g��DK��d�I��c�N�v^�4�f�w��1O����1>��  7B�MdTS�����q����U{�-1��U���#�ז��G�睁�k���?��*�����їb�o��)��t��<ޖo�@��w�X�ާ��s~�{����҅���gh�X,U�4Pv�ܔ��J�|j�"�9i�.������ӧ�����r�}R������,l��'�-j����!-�§���-�ޯ�޷�y����"�C)3N� :�W�$�T�����3���B�)I\��^�� 0��x-g~!��q�[�2��D�u�1z~ǻr�C���}>�~�̠-c?E�#k��F��^d�!���U3���Ue�]������Aj�g���mȠݠ�����ε��r=][Dn"�Y&����(���4�?�nw,��+!u���Z�-�b�ڊ�[� ��-㘸A��ė��U;�	�����6��U�����z̗�Q��ю�|IB��/{Yɞ�4_u�Ms�a&թ��ҟo�^r�uZ�4$����I���0|��1ޥeE���ij�{����
C��$��|���H(N=���<��i��࣐p�+v:~�v�ڿ-%F��S�QNج}j��E�d��`Q���#��@�ϾD|	�M5�I�Mi�-�\nYU���+�U�/��x����l�1�*<2�/����8`y�s�̻ �E,�ZC���
�����&�7���[�e8�>�Ӽ4G�R��d�p�X�b�tfg�O!V��D�O;Jc`�'�k|��(=(=�W]���V�N�X`��v��V���� "cAyo��l�*Ne�M?�bCP�\[V`�n�z:\E{m�V��2�|�>1VH�m1�Q�$��Q�\4?�Xdh�vB�M�IO�f�>�'���ѐ��\hj�e���R�H����Y����Ęg{�*�\O},͸_؟,���=C�w�C�|��*�f��މ����4�*Tō���y"!���)|&��(��u[&R�>�^�8���w�-����}�rkv�|"8�[F���P�'��j������ю�=��O= w����$���L��hP}�5��OS6Y��+-�W��]���~kⰫn�_?ܣ���4�E�����r1	��
�4)ղ0%X��,�[0�AN�V��@�jY�/��fّ�(ݦ���(q�����9 aI�s���mu4���P��:z>ǝ6���1�zteOR���<s�hc8�zuw2�h�8jx��X?s�M�Y�ሑ�C�Ow�H �Qq������ɵ|��c1��y���eǋ1|ٓ���}�2J'��G��)k�:E��d�\.����G�B��BO?.�:������?xMY��g�O��rM�~���ۻvƹRvk)��d�"x��.]<C���&I�|3�W��r�˻�|A�Jm�XA�m�r���^~e��	:.���-./�<�\��i:� |�3����[�~��ф���5�>h��୯[�وz���g�}��w]u����֏֯^��
{ޝ�_�[|���:ud�k�G�uX� ����4�<o�~�fy���B��� ��;�l�����~
�l�GP"�	�Ld�kͤ��O�+sBF�U���kb�*�+U`3�-ޅ��@��w���9s/ʂ=��Ь�>��`JU�Q�V��Hp���&��s�$R4(bFǑ�H���@QY�I;�a0#�U�*P/}��l��j߷h����7�I���ޛ�d��xz�6ū�R��w�.����}��qMm�hK������q}4�A��ȉ�~� }��҅�*�i��,�K�'C��} Bf����^ѷ��rB�w�p7}q,���\�B8� �Oo'�$�!�{{�nH�ʐ*p�k�C6[��gC�u��T�i��� ?��q��>r�Q���{{�ҩJ�d��M������uU������@zW~�8��wX�[}����*?K?Qm�gp�$�k�o��v�����&u�X��-}m߫�m����Q����}f��Y�h&��ίz�:�
�/._��/�D�����i.���l�1���o��/q����:�7���O��T�a�0ؗz���<U��v*�w	���o��%�J���d��k*[�eO�8��*���*Z���-�@����q��g���t8.՛�8��Q�0��,�{ҙ��Ԃ=�v[\I�RR�n'�gv�ɥ���t�M�;�Q'� u����
{�o����P��躏o`�C�<�T[�noq�tFn���B��\�
��oAR6Uq���7CЕ�ͼ�+�)gD�K\g��6ۖl.�L�˲�EA�e�q�fϠ>ێH^
�D�曩ϋ��^G���ۍ��5P2���j��A?5jqի+e.�!F���m���H�Z\Sm�A(�e4�??S�~�l�YM���ʷ9k��}.@ӏ7��◥�>;C�A��ly�y�FY�宾�P���SS����L�@���3��f_�/�ЧKh�������iK��E���]Y�V��#={�E��]��e���3�
�	����F��6n�i������_f�����O�vc�Z<���MF���o�^�?|w�:
'��F����iU�\_���$N7x��*i^�Z�����5���/�>�}τW�QmҼ�:#Hw��<|9���}렑�+�k^P��g��	�tҽ�]?6��[�y�*F�=�D-���8��UA���7��_=
yw����lN�n�ԅ1��]2�o�4��bn'5�Q�X�����e���~�9���>X�-�Ǖ����[k�߻�,�er}�O��Q`���Ϗe���3�)�	�^��Qs�~ՙ˯�?֭a!nܪ�j�Q-+1����ۘ0\Lm&4�EP�nk���>���h��������m�A�AW��K���.��ݩ�����Ó�_^�ܾ��y��ɜ�%�A�v(��s���4�UiL[�A��a���X�6_�B�~��L�9�*��O(��c�/��#�F�H��*��bMg���n~��T�~����&��T#�U�0H8�n���s��`uҰ���D%A��E����)u�
L����B�hw9#�4��xa�i��"��B
R�tah.���j_ew\�8�N&�������p$$c��������0�k���YI�&C�N&'j3C��'�nD�4��*»jM8R���ޤ�p�Rg%��{�5̣��Zڧy#��ͻƢ��r�w����f��	��P�S�����Nhwڏ�vUF�p��ǜ��a��*Y%F8.�e:E�8܉�W�{U�ϑ���ф���?����M�n�:����g�;l �P�6�5�� @�Cb�C��.���v���$d�tw~:��r��x��[v���߭�S�oşZHoOOO�T�zR ������C|.�G�v8c��D��q�+��d�$�e��D`-!�L�8n0P��31r��Gd�G.2�V
W�a&���%�{��l��Άe�	�tZ��1�2^���(��� �xO�y��z\Ap����Q�%&����PdW�����!.��<1����=�Vsd�%
��_.���qΝ)�7�w����{���;J�a�l�=�l�i3��+��+gm��%��h�q
���Fg�x䊅ն˴i����9�����m[FU$C�,s��p�g���g�k:��f�����tL���.�g���CNr�ǂˎ��?��(!�Y?*����Z�ɢ�n����N8$���r]��.��>�6�Q�Yts�}s���N�l�wɶ0:�ފ6��.�.���Zs��_�_�*fGK�zaD��z�ى�тI��JQp+���tt�jkj�N�����4��!��T��if�Y>������[��[ �Ϟ:���+,�w����RVҘ�)�� K��=��M��5��n���F�]QNb�ks1|�H����x�,��.��.EQ&�/0���Ĺ>(Q�B��9�*?��
K�����~�'�"������ "1Ȫ*u�M�K~r.y}���q7�&.����'���'S�	T@32�M(ᙁ��J�R����ə�6�m�i'��f+	�=Q#Ǒ�8���7Zѣ���X-��^�ȔGzc�����'���������US�c2���^�Q�Ͼ���Lt.Bw�~E�%�o2u�?�;�OC�OW�J�A�o���A!TQ��GXY�`6�g	��	{�V}ta���0�W������l�����l9�O�d��d����=���O��9>ac��P����-뜚4�ѮH�<��.]��#F�&ּ��+�Ri�KQ�e�b�tOK������=�o�����b5.�� ��[D~�*U��F���A���c˗�6KyQ��'��to;��>O^�\]�r�P^EN���Uky'�5�ڽ䓍�v��^Ζ��<F�F�V�|!�=[��F���<�Y�bO¨3��eG�����-/Q�w�]���U�M�����%� !1�������FUϗ��̄��\߻P߻�ק�W�Q���U$��ޓ��Zd�������& 	U�/�UM����l�;�����ֳ`��T���J~c�q�~���L�yƢ	�!�
#���%f�B#̆��I�{8�pLA��d��A��2��ͧf�L�C��]F��O�̉�=mMWV<#��:�U} 6^rP����p�9஧g�G:;<�fX"#���^g��}Ѳ2��,gHP4�-y��`����.ڠlē,��g�Vְ�hGy�Қ�f�ha�w��8I�Y�;�?��d;H�Q�3:��9��4�/����S������AMA�Td�Y�:��^���Q-��N����l7䵌�c�����)���!f�պPBH�d��<L�F�E��tq*g�He��$z�e�YO`���O<���:���F'�A6+���&��~���ĝ�*G�b��|���jҀ%�B��'w g�O=���}��Q�q��b�7�h������cE��Lև89(�i1��?�02���[�.G�{
�ݎ����O^�طg�ZMТ�ŦAU�L���X�ےH2�2}���x��ˍs��\ԴG�3����#������*����b�Gr��8�qo���+S�̹|��h��*| ��np���������k绳�|z���`�I̜7Zz��-T������G�U.���:�����V��g�K�#O$={����͍���G�M��c�H1I827#ߘBؘ��gxe��t��(�,��ɀp�A�S&6�����I���H��g�ɪL@�ZرJ�Z�`����N�P�Q�&�CB���8|�j2z�jz�j񒻿�cB/�K�m5mGr]�Dk#�ʈ|�W��]K.ؗ
B�$�"X���ŷ�b㶓��GG'Fu�����K��'�I��D�lY��Z����u�G8 �L{��7��9l��Ȥ��T�d�J��B����~f��<М$O\�Z�&��G^�$:��ڋ`�����u�=u��s�Ou%u<���9�ٜa5;.i3�4)��P2����,��c��k�����ۃa��{P�����IaS�=��޸�;��W�
ny����V�,w��8���EG����h|����K�Rxt�-�[ca�QR	i��{݇���[uO����0ț܉��?Z)��q�o����Fd��㢽����Q��j��x1�{���u�p�`�sc�[$�����iP_N��,�S�[���ï1b13���C��6/���ɐ8g4-���a�B��|�ޔ�f�q�f�<�7��mF'���Ws��4˩�?��y�rξ����a�����u_"|Po-�T��2�@Dg�ə�]��(�N�u/�o�)��"���o�6E$鿈�X+�Y��F��%^�΃�~K�1��f�4h�va�o����}z���-�w%�����;z��Ho���ᄍ/��ŀ�:��u���N#��]cB=x.U�^�F�:�:��վ��ɜ���ǣ��k\X���7�dT�uQ���z��s�6&����끳ӼMЎQ�OEG�zsL��k����vT\�  �u�+V���T-{�A�z�%����"�b���\�����ow.���c_��Y�f�t�D�`���.~�F/fJ�0�X�f��� i�b��:D�6�l�=�'&P�F��Q�*�M����ێV�酆���9>��<w+����>�;͆垙F�ӱ3�7.�99U�):��6�aa<�d��(�Sp�Ȣ#�[C���ޱ0G�4y�#�y����G�#��*���=㢰�����~X�gx�	:+[]~z�"\u������7�y����5�)8wH���b��W:P���׻^�y������͏,��!��0<���qw�bk{<��lze>���	G�a]Bǌ�
�z����WR����	���LlU{͏Uc�ڶ	ת����c�0��W����IŨ��Y��4���֩�:Z8�<�̽�E��᳊�C�KAS\��?�Ǻ�~����S�To���ZcS3aɉ����ū��	w�O�G��j����+���N j�M��Y�|<ݫ���B�4��	쩱-�
�N�p�r�^S�8R?+t-(�1�N稆-N��x�]VR�"�x�,�bG�"(X��jq��n��
,)�b!.wl�����O>��X�B�M;��<�a���+R�׺_Z�MK��	��hg�|To�UY12��V"�q+��\�/W|��l���~CD��GU�y?Y�/��<}���BH������{2m������4h^�PMl&Ycv]����i��� �h���N�l<l����^8���2]�n��I��^ۊ�]}3�Qh_������KL����u�aޘ���17<�ӽ�Z�m��et��o^|λ�V�˛�'�}t֔�zo�	M���3����/�c���i9,2�6�Y1������9M��P���Z�;�%�N���^ⳕZ�5!P3�;[�ǝ[p}�9�aE���0`�C�-��ڱ�P�!*~�2٥8��]/�.�ڝ���r.Ή(&aĪ�2�-���`"c��EɿV�	?BЮǖ���$b�����͉���7������Z�'>�a�� @�?M�Xg��nQ�w}��8]��̊4����cO/(�4]��5��G����A�H٪h����I�bfb�4���(魫~�T'�[+RJe|����,����+�����]��B0�����=*�n7��5��O!=і��i몈v�s��J�ꕄ�#j���:�_u����i~�w���k8�Q�`��ӄ�řI�SS�����^
3Q/y*��[��'��%T��p�y�FK�V����˥���e�N ���� �B���%��~n�����2��9t�
��B�~,��K�v�.��of)�]��	�'�C���Uj8��1')U�Vn�9�[����=_e����;��J����T�U��Wض��V�u��ηN��Ve�îL�,������R뮍��u�A�;�=��m61�x�7Vk�[���@��{��B��26���X��wnc�f��y��%�I`t�ʘY�� +`���p�4GɅ�Rp�A�P��2k��c�"�>��[�и����^$ޛ�pzd$���� @U f�,7=��0?���1JM�Jn`f��gLF����,A���'A�C�3���o����فEQFGg}9���_��W~�'��!���c���|g�|G-�0Q����M����ⱟh��������M�f�B��~����)bW��]���J0u�},�E[A��_�N���֙/�Q��"�)����ţ���K$�J�a�/I}f�ɤ�a��w����z��ik���Vqo�*��qd�n��z�T�GE�J�� l��^�D�	=y	P���>K�R��%��R���{��<b:tĻ����suQO�H����me�ؐ���\�v��/�M��Y�d�������/�ο�m�[��Mػ���������0/�f�&%���T��9����	D.�c�ψS�/4�l����2���.Q!�I�)�d{�Ay�=97����\[�BZۗF�j��^أ2��)������Ͷ�d.�G&İ��ʮ��_w����=)���X�Y>2�<��~�&�KD�,'H+�8�Vt^,<�GkCJ�QR��W�d�)Ċ�17,�4c�B5��
*^�ʠ��P��ί�������&�SK�̇��뢸 ު!�}F��JG�q}Y?�n�gD+�?����h5}�%����1)�3~t���~��މ�ohR��欂�Z����<�Lˢ���^L:��91���#�G-o#���l̙��6'!���n$,-��Ȱ�Z��F�EGI�(�j^��䉯?"tIbF��tD�<��PUY���Iz�~a���������D��p��)c�w$��e�q^D��M�w�/�)���;�w�}���J*Y�(�`�v�b'��~,��;i
m��m�'o�h�~�Iא�\�/�܇�p��=��;���.o��r`}ĉn��8k ]�#�|KA�i��iU�$�On{H#�"�l�M!�` Er�Px6}M8��$뿕�|��hÕ�3�76��Ǔf����>�Dtp�蘴�=��h��]G�9�R��<�ϻ���k�#�.���F��)��̓/`e����ȏM��2\"6�2t�`�6������.��
;��\�wa���C�A�~[B�D�9I^�S<��|��'Mj�ܱ�r0�̃%?����KI_�7�$%��3'��i.��3���<�X������V���*��K[���ʯ�M�������s�Xӝ>�!�ә`���6[T�F��(��m�D9���|h�i?��JC'TR��ږ��M:��h���[�'8����d#~�Cݍ��^E�ş篳������]������uY��%��؋�G���JVOP����G�]ڊ�ep>�|4!���$=�%�(r����3�0;(�Ә����\emtܧ��Yն`4)_����O��]��%��H�*%z�'WO/ B�,�y�����Ю�RT]����qE�w���(�6�������R>7`+}nt����ZT��?�{��е~k 2H�G�֓�Z�gG��wIތ��e��;s%Js�f��"�Yh�r-�S�0���'S��R̉��.B@�a�s�a%�ք�J3�0��(�U_�>mϷ���Q�r֔��5���W@*d���[?�:,��M�,��")��JL>�P�S�B���:i�gIK͸�Z��#�MNy�8����As�����@hj0�oh;�`�"������A��PqcJ�d#Ip���~u`�``���'�AM�%٨#�وۃ�d21��ʡ[��ES�?T���=8}~����)#[J�W���{Z_����."2 +#Q
����6IGI�Y�"*Җ��g4pt�:�}g|�<�F�t:"����@�Q�hs*��T�����������|�X�qx��L��Sg��w����+���f��9� I2�x7�Ĝb�}���Q�sh3��/�[���g������-��û�fa�����/:+�hW���0��#0A>�͕�����-��y
�gd�\�,�4�]�%��C8�6��9Q�2���O�%��u�-�����l��D\��(F2�>e#*�3���h6�^��v�y��θ�ˮ��-���9ֲV��f�j�r�8�޽3 �3Ua��Q+��Qm����7��+H]CCn��1!S�vY�w�g<�W&G�Q�c��&�&䘃���h��!�<�o�e���h'x�U+�&�9�>�^/��E�k!��oi+�B� �/Z@�F>�I7�Sf�C?���Y�6�������HI�/E���b �b�b1�)kDË�=���{m��U`����Ӹ��������f�(��I�(<�,C�
�/�g���V�������R������K֨�˥�Em������!�%�ZX��PЧ7��f~��9��y�h�X��eT)�J��?Hp`��r�sm�ERŵDp��4cp|%$K ���)_�yv�!�|Ì;C�����:nծp$��^#�Ms%���
��	�����K�z��((K���T�^*$W�✴����zn��ض66:�}�TOk��l��Hl�1_�5-��m����F�1��β���r��b���Q��B�_?N�MkPM|Z~���!���M�A��$x3k;�n��1{���#���9�~ �<s��3gh�(^D���4	�kf�$�#L�w����cM���U*y���o��z��} ��JJNƶ��}9�~=k��_&E^/E^_��h����worZ�{2'=>V0Q����w=Y��O�ޟB_����ǻ���7����EPs��-�!�������2}h�l[ |��[ˈ�Z2ѓ���"I�Ѝ��SD�Z����� �]���l֎�����b!*�С��3���>')q��������E��~p��2��H�����v�?�|4M�<�YM:�m�rwT�)\�k����zAT�����ME���S���&l���I�x������] �`ަolX�4ؔ%�<����6q�%5ُ�������kq͈ԭ~eH�D�X~�0�(w��?�*�>3D���ُ��i�{���f��g
�>��>�dߧf�C�����
hc�cu.�?`�+�����:�ѱ�WN�W^�����̳��<�\	����U;�gB�4If 2�%�<��m`������oKB��C�-:�9����d��
�h��τ��M�G2kk���r�T��z@x�`x6�V���짭Q߇�엟;u�|.Gĳ�8��S9����zX�{���T8����x���W���� {P�`W�?��v���z��� |�]���d�2�_��U�D,||��/T��q��$������� �� cCV��M0�� �~���t#���	t�о�W��:���Yg��%GNm�~��3��AffrP��<�����C^�zE^�eb���e|�d�����H�(a��s� �y��i>"����ғ�E��oc��x�o�|�p���J4wy0�GⅪK�aǢ��
J� ٦)���,	xP,��QP�\b�n�ߧ��
4��T	&M��q�h�j{���wE��Rv�,��;"~;�OJ-L�ur݀��8VBP�>��+���<^=����۷�/�Ї���ǥ]��x(��^��B��N0�����/O�v��L5�4�w0]��#s�}\'F[����r~���YO�[�i.d�%�-�cyCO{���1�X&��(먪oeo
9
<M�Բ+�����b��?��{�D�\����`�`ψf{	�O��׹��Q��?�'_T��Ղ�W}>nz=9}9y�M�����=ۂ�_�}}����GC�ƅ��C%N�_5i7�_���0vҤ��p)�F,k�*� ��2���׿���!��D\���/zH[�
�<$9�O����4��@��B�1�i"y�\� 5:c?�/"0"n+��"J.�#q�^S_(���q�W�\�o�1��%D�F���b�,�|�z�	l�,k:y(�ylB���ݕ�>�����.���j�P�#�y&X�G�2l*}�+|�T����GEz�`�l���j�]7�7~�b5�S�\�4Tg�ձ����ڑ��%��m��L�݂�	�a��{�GL��Ϣ"q�A��ts�-� ���32W��0~B������?���uw�N������`zuT=
�Ne��J}Na��:Ą�;�H��꟭Z=�@%I�؊r���JƗk����5�_�"_>y�L�hZ ��
��c���qj3�6����l_[[[���_��q��@�~���O��Mlg&�7f��	���x�㹢����_DtJ��n9^O[0H,A�����9c�l�L9�Q���S�E���#O�\=���_l��t�w��u�G�``BO��:��ٞ7ω9��zg]9 �d��===_�d��2�I>���ݳ���m �ͺP�l<FW
��G���'sa��,��E��&��E���;����xT��@��Mb��R�iow�	ݻ�u٢j����������d_����y&�U��L�0�d��,��x�Ç}!���`"w�����I��|��d��8�{v�Ƭ���u9l����,�O�RF��p1�&�,�G�F\��d�\t�W�<�",�!�^�/���,J�E�Q�<��5`�#s}Cݘ�p0��[�{��?d^�x۴i������`���N��}>ɰ�a #uE����8o1�b=M4�P����t/�I�>��A������ �@�0U��r6y����Y7df<~|��>T����m�|��FAΙu�Z-�;����I�l���6����Tn��cB;Z#���A6Š����@;�+�\�s<�Eǳ�b�=ɡ)�K�˛`�N�6+"���`��G����.��!��!qa|7{��Y�-㺜������sf�|/ѷ�p����:�����.�ƜU�{�@����$O�ְ�IsNr����4͓�xXћB��(Ǭ6�̚�<C\y�n�7�'��B��׺�1����Ź �3wƱ˥�u��|��Egzś�(�@s�S��i��m�F�/gv��"�����n�_5��-�:�鯫�8wnt�>�o�)�R�U�㈗�ΘF8�D�OW(8��1�(n�
��Bs`]��T8�����(�:ŚA\<�Z���uTAܲ�@c�q����+8�Z����NQ��Rw�ْ>�^��R�_tPWW���O�+;ul����Qe��tO��?�6�|��y��ȴ}ݜ����t���]p���-�w���*'�д'�Č�n��iT+���~�[2�1���o��i�wOj%A�<�cu =!���~$MA�	���;�(�������I�a���w/)ˮ���.?�:�
�����͎��4�oW풾�2<c=+Z>/��j��i�<���~=AJRW�V�Rn�z��D=����/K���f����Q�a��i���a�HB9��{�qP��Lm9�d�Û��Mg��#����{V�m�I�~�@�I���gC�B�(�.�GM�5�T
�]� ���I��x3}���]����z(:%��1܂�������E�煶�6���A�$M�s�=�����T�z�ޞCk�T�M纟� N7�̥
���0N7�::F1#B- �a'�� �o� @�4l�NGLY��3}b2�:rH��!a�*�/��a��#�7f�u)�E3X!?^�`�(6d�iE��J8���)}�L�tf@Ϯ��W5�f٩z=�@핃M_��I����Fg��k��.V�΀�7��NO�)�D�4��� 0p������C�@<]�`0������r�J�IO�j��fEp;S�f>��ט���|�oZH#ڟ��,	����x��a�j�ث�G�i��/@v�ꭕ�E������Hi%������'�vRs`:X��b��k����t��>�la�H"���������\�oն����E����}�t����#�|�p���qY'-r�z��_оv�2|>���d[0%�u�G���0��Z�^C�X�\"��i����*i;��b��mz'+~������&�̦NZ��2��������ՇǢ&�Q�Ed ���X=��i�����V�E@"���cxa����-�Ų	�I�f�z�u�2%�S�~D������1��Q����Oװ��`��+N8ͨͰ|��U��F��h�/L}L��ŵd}�&(��.Tp����cNT��ǝV�HK�����疵�1jO��ts%S�JO�rAZjvH��C�Ĝ��3ׇhMtٮ@s,bj���Nv������[�*����䑪��GmA�$�Y^���R:t;���I�T� _�hK��]��t"�LxZV�v��!W����x���Ê���\��g�K֥;b�=�(��T�O�o�-�S�l��s<�g];�����e;"��[��ؤ����;��g7p���bۛs�/�/�̛��Q,qJ_�[�V���-�y����f/V2�_��t6�ۄ����{�x��|/�HNeOճ��)��|>��-xP��ܲ�(v�\�nA��}{�O�Ck����m�
���d�~#���[�ж��d���]�!V���m	,�Xw��T�����L�u3����b�I���2�v�,��8\��γp�9Zߢ�aWr�=��	�t�G��g�q�[��^=E��[0Ŧ�c�Ꮜw:��eC�v���I�b<6�O�>�s]�BweJ���O�x�#a�5��lu��r�(�få�4I�y��C�}5��>b���.d�i�w�G�@ Jқ��ot]R&�t`��T��Lu�t��Cp��G �j�&�]��26ڧ�$��ns�`�^�L�Dxq��{�Me��H��6�-QMJ�fkKy�����4��v%�fh���������+ius~���o��tf��g���e4����[�3ժ��`�GKS��j��|����5 ��N��j�FċI��H�.�7�[�m�����Ü2��Eǝ��B[*��g��gxO��
k��$'�$�� ����^�B�Z�1��gf}�vb��8E��ã��5K�~�EO�oݰL��n����a��5@ʿS�A�g��MIj��#O3I�we¦*���o3�I��n���9_��*B�0@�6�@���S`*	^JVkQ�I9Th����f<�z]ڴ��EM���{@����/=�=&� B�9=���.m��oa�䚞C�z�B3"� 3��8�T �1��?�hX%�*�/:�P�y�'k����S��	������	�@)n�& YΚ�0�]`&ǳV��9/���%lWP*XO�ʟ#���>a�a�%�6eE���J�U?d[���������r"䅳��Ԏ'x�)ro��1R��:��nJ�Q����;���㥨"�#Y���{n��<a��zs;�+����޲v���:�W�����ؗ�$e������70�;Ǽ�K�A�pA7�$�S��s��56eo��m�8�ĶH�x���8I�-W�� d�A<�+�F����\D[4��L�%�%�fJ@$�ʤ�������.�OEf���)�yŬmy�o�,qA�u�sG\J[?�z�[��"��i�����P][*�<���
kRK���ayR9�s���=[���RE\��7"��צMx�&�3	�u=�U����&-t�&W̛Y�Ux��&�E8��z�L9i��;���scL�M0f���ԯk���IR�����c��	藢,�������'n�.jn��0�Y��r��1����5�?��q��1E�
`�h "k�׹��n�N�~Q?��jz�&訩�������TJY&�pa�`^�߃k�A�3�>r�:a��~��h�rUiIo�1>�L�n.$�]K�TM�ga@�T�m�h����} �栉K��Av-6�3H��$�N��#�t@��	0$��3*�
�Hc�v����!���j��Y_��j@�m}��!+�����lc�ǔ%_W�0����J�����FRi		���:�~�~*�;����a��h�K�`�I�	��80^��DQ����$�O�<��Ӂe����®sH+CPѻ��]��aJ❩F�Dy&�&x�/\��](Kl��Ǒ%�]ts2�͉��|r֥>%Ӷ�ƨ�:���)olG&X��$�t,�u	�i�B�I�e�~�W��̐cP�A������ˎO׀�2�G����1V\��J&XF�cL�i@�S�h�̦�[5��BF�r�(4�6�+�J�k�=g<w�������B?H}t_#�,r&I<7&���
�ݕ_��e�?;=�ݜ�˖w�=&fIM�����1_C�C�Tݭ�wi�O�m��s�6��t�ҀX�s����g/�� v�����&��R&0�:�*c� �ׇ>do-HMͥ��MQ�v�F)\UI��&��sTV������p	d�q����&�%�<+�hi���kl*��1O*-1,�JO'6�DJ�f���J�AVΛ�a���=S���'&��#λ�@ -ב�$� 3�Fa��^�	��e�ˉS7$}���i��c>�D�S�M���0�ݛuhb�o�%���Pcn#5��w���o>�9������).�2\p�]�b�a��ßdFe(7֢��b�h�އ�J��Q�'LY}D���7SS��Ō�O������٘�j�X�eL����/��hw�&�"�%!m��wk���oC3�L3����6`��AT����K�lytT�G͌������A��Bf]� 	D�V�2ٍ��{�?Xi��c�]���Z��+]O[č?L��3��l1���LD{k�|�8w�jx�������ᢎ�7+���P�g���1�>����B�CDuJ�w̾;!!bYn4��I��r�k���������M��>`��k�j�r 5 ����I �M���UA��)+T�!� h�d�8�=��-h���=�O�S>�
)#	��?�ݘnM���_0U^t�L�o.��G��6�yf"i�>����\�$�l}�yTh��}& ��d@(0���7I���x͟gV���a�P"Ð�]6�f-�!b=����h����<?`��v�b�d�Ĳ�60����48 O��bX�U��Q�yl���~r�ʖ΀&w���b<����0���i�y�]�U�#lo��GM˃�*XA��(#��4!\5�� c"�m�b�p��Fq36ޅ����]�_����)�����E��nU��g����eb�!�kŅ�>z���4�?��D��k�9�{�oW��>ľf�u����f�����a��}�+߳Ta�b�5NFHb~�-< �z�V����!&�v��mLYT�M�n�QQJ���0�:!a����$��P�&�?� _6U��dl231X`�|���&vrC�QZ�s���z@�#��͝��cdlX1���b2����*��r?@�m�7��zֳ6�G�w=����q��1��w�����g��>Jo�D��w���3`h~��W_���R�(I>��^���u3 ���J�����QPza˰~�����i%�S���PQ�Mx�e�f�ђ��
�K�i	��t���:�(���D3S�*�#��׾}&��A�fUȁ$]~*T���j_���	�a[`���o�Fk�|!@���5u��Dȶ��UGH���ԅ/�|����2e��\Z��v6��C���1 ���Rn�`*3am(�<�X.3��1Ut��>Jt;'&$�U��ғ0�+�����cv��Qv���hY�#f�DS2��Ha	L���h@24�2v�dsK�˘���:#!AL@�T��GM�{vi��Z�=al�e@�9]I닢ʚ�������P�-�m�=&fdW_��W�ΚL�:΋�;����G�	�<�N��������}�@t��2z~?2�/��vmCO��vu�mN6��Č���+�����)�,e�CLY>X���f�@�Y�W���K��f�.Ώ�������ĳnv�F�����Yw�[�[;}TԌ�1��^X�c�Q ���cW0�����*��[��Nd{���f۴�٤m ��Mc�����h�����Źw�ZnU��v�lM�ڏ%$0p�Q�ڙc�	.rv�#�ԙ;X����� �h�X��F�8���l�k� �KO���"j>\>CåqJ�"	4�lvH�b��_��s��/�Zgxi�|� :!_bo�����g���>�|��,�1��|#�޿eT~C�ߟg�2:�#���/ˌgʙ�����u��g@����笘�Ș��M��]�t�mlM����N�L��ޱ�	LX$j��:$'��z�>(lT��
JA�ǚ7�}1f�z��ly�ߊ��1�qz�olm���E��ں��]��yo���%�� !&�M����$[|�Ж��ڲ�����9���;k[��Q�"�ykt�������%��Vc�S�g�,����rXA�P88�������D�)j!6L�D�Q3=d[����aV(�.@ ��T�,���!���&��YO�-��H�9�)�=�F�d
%g0A��*e�i1�IV��Hط���Z�7%
�F���l̀��Dː�cGO��|q�?F�!�)P@�l?���_^,��%�%�U���'�6/FP~l��-���DD�m�~.���{"�th40W
$�y.�<��>�A5
���Q獡IMe2dx"4���	+%U��MAS���I�tG4R�g@@#3��d�խE�M�(m��Cs�.!������,���]� �1\��~VO�ct����i�A8�Tf)�b�ͺ�Y8�4��B1fko���p�2�����,��T3Hc
ʆC��?��{��] �};� �`�]�����"߹0���	J*Tyy���@&h��M�	i�U~#��b:Sd3ϛ�	��x��Sn5��� ���\� H� Mr!�`�2�ߋ.h��
+4SR��C@�AI�&�9m�7J��g�️]�,M�u�ZA�D��l$�V�.%J8����!~����m�.�'�Me8ԛ�-^ԛ��c�d�b����W����8$v���|!���M)pr���Q�b�!�ݑ��Hd$�I9'y�@_�����˚�y�Qx>0 �r��c��u�HE�
߿�E��ktB'S��6I	���4x_Ġ4����}6��R�0 ���ޭ�e7���`�h�&�H����`��[�y߄y� 92J�!R�2!֞�r��]٦�ϰ�a�����)ۼ~�=��b��=�{d���(��|4��s�&k�a��w��~�~�����7v���ܐ(�@�M��#M�1�Np`�V�	�����E3�|��Y���bD�4(������D�֯�,�[k��
�%H6�5���h=�Z|����_���g����3g_A!���+�ב����[:������;O�ŮLAH�an��	��r���9}'�2'0ڇ7�`���n*q�,,��(���)���Nؗ�(IZ�*ӷ5��������Ylqi��V���n~*'�'p�ђ&C5fp�&�9VK?ʓ����1�	��g�b��>�Hc�9m�	P���[�U>��X�=`�Q��0��u�)�H�($��YYp��C����	'�zx=
d�#<�fP`�Hkz��	��U��v&�>_��&붻o�ࢃ
����@�p��x`�7	�F�Q�Y�O��� �@́�"�	���K��䀑��X	��6�>+�����*+՚��%;y�)v��	����ο�{饳L�16X;ώ6��Kl,4-1����S��ؘ���\�Ё�2ۃ�jl�)�m��ocs�_o�P(�Ƃ�D��i�|���|!����粿����	C>a%7Z�L�A'��������Cv��U����=��9����عW_e���e_}=@TR�Kt����&�luqU�m�g�E�T�bJ���a�"^�67%N�/��x��f@ln����[L�I��2��a�c]^lw�O�fF�L��e��T	��̱�R����p23�a7����͝��\�tִ6	�b��H�w��-6-�|{&V/��#���$3V"����zT�|������H��,����@��(�L�P��3�ϸ�}1e�
J�go�l�Y�q �D�����{<�m&j|l��_ؤ���$6�ð��ČBӕ���,�I��<��Day�Ċu�E	T�o(�I�\޸�{sËƲ4D��(�����?�؏���$�4�~�[[!$�d��4s�O�Us��Y 1��+�2��^��.b��7�3�z���رJ��>.�7�����j���wG���/H�:�<6@fZ�-�gV$�5a���;�Μ9����w�����}��W�_��_��_��?�4��W������� $�`��(�Ŷ�����2�?�\�e@����Sz>Zd�'�6�n�j~//��L�U35Q?�ݔ��L�ϖ��`@��h�ZZ�4��1=X��t�� ��IB�l�8�>��������s��/h�n�������w�����+���/�/�?�67�5#��x
[`�h�!���mq�����`h�K����ED4	3�� B}�vQa�Y�2����&���콚W���S7/���8�)��`���		3�rP�_PC�GU�w�Bpg�Q��2�ى|͡0+���q��B�p�-�ѳ�_=Q���	��n�t8 ���L�zkB~��l�[��d��� �~��Ә�+�]0Qe�oA9�$����N�o6ѭ(��/�\�"&߇������Dx���Y����Z�7��27�m߄G����!'1؊&*ˉ.�t�]�`},'�|2�X�l�u���:����f���P��w��JMZ��I~�ۏ�+�`'O�Db̌��1*�͒��=��_YYF�����o��d�Ʒ �r��a�{����4	`c�Pe��՚]Z����������v4��燹�x���P�o6S��d�����f���`��I�܎]�p�]Ԍ���&2d<x?{��K������r���{�dg_x�]�vYO�Ua�4Ӳ����Ul<� �K9M�t����'g��8�#���|�^c8v��8�{	��Fǩ��Pfs.�Mp�5V�v'�&3�� {���M�(NӦ�x>�|Kn%�P�}#��Ө��]���Y�����b��G��2�b6Ll�#zg�/a#�th`��B���̭�@0����ɚ�Lu3y�#x=��w�k��[Dq�ۜ�(C ��`	�픹9�J��D��:mb����:q��)a$��)�ݕVb?�n�|$�]��`���a�|����闾�e����]�|�]�~�mn���+��ٳ��ty̶�Ƃ@�>�9;th��,����xZ1 �WD�;����ߜL����aN%�v+�%�}�+s�l`/���2�![Z^B&5 �7�2��4>S�pmjf#K�*��B���1X�������#��c�������s���-���s�y�)�~�*[�\cSd��e��-�K��D-�2f�`=3/bռa��rKA�h<ЫuE3�C�|��!޳@�շ-�5��+�cPz��F�9w�,1s�W��y6<'y�D��DQ��������W����U̞C����7���%�h�ߝB�@��.<S����
m���s._�er�tCL�W\��Q�&�(,�{�M m���B�HD�߆������e���O�W�;a�r#)'_8���B��Y҄�}���~�����:u�����#�ԧ>�.^�h��j&��B��&�)��P� h�������ǁu�	�.1�,0?������W�������y�2�W�lD��M�����ሕ����2p��֒4  ��2�֠�E����¢a��SԂ�6����n\�fe"�M��|�{�%���F35��S��d�Nc�^d��L�� �pK3n<[ĈZE>@�'�Ӈ�33��$�0 ��+�~]����(�v��<��w*/HW<}4�.�ܽ�j#gzval��Ā$�<�P�� ���-Tj6���e7΁�H7�	�!'3�����{�!}�.��r"����@��[!�~�<N<�CP�˻�`Ep�&(�!𥪘�@�l?"���{�\D0N��m�3�w]�ӽ��WG��T/��5�31c���ba2�w? �����q�@�F�6F�v�s�A��@;��ȑ򥎆yw�y��kc�c�0�y���7}�4�!y6d�K,x��မ�N멯�L�UveM���_Z�y�J{Z�ai�G�%�3ʫM���5a=e/��{���aW�]Є�y���K���/��#�F�`� �X)�$˄��F,�{����̚p�5)�Dl0S�A��@�W&X����6&YhbUJǬ�f5��1�L����H��oI�~Y�]͖i2g ����	
eJ�Z��An|T����M�����_���LŖ�����o���G��&����7�h!c[8��P`xІ��&�R�B�{f��kx��?0�Wnj[�Б4 �N}�}s������$w=�؀��A�pFh�:n}6J�D<_ _�1K�<�vw����9i����B�n��w��v{=�%t�k����w�Җ$��Ow�<�L �r���Ӿ����#�I�%���f�&�41�曯�o|�����0 H��v��p���l.��b�j"4��;ys�v�ע 8Ω������o �WWU���d��l�s�6&W������ҙ�ahg
d��@�Pcؐɘjf�[gr˸dƏ4`��01���I��Q�8�K��9?�WE��CL`p@s��4Bs���Dm�]g��ZKɖW�Y�8dW��3,�-C�2drh��d��R��"$$!!!!!�ve0G4E��)�讀�����w���PS#^N4�������lz�U��w�D����;v��X�\G�%�� ��+�t��IS�d���`^��[�!hJ@J�П$ʣ�a1*<�t�C5��UnBz�f�s^���?S.�m�P�\���L��1�:.��Ąkl�Q���0 9�6�0n��v�D˲�� *D~S�66�����c���6�ٷ��[\^F�7`|�^hF8-��|>S��!1 ��q�Dl�!�1�@�~$�~094�,d�R����m��MQf��Sb�Z���+"��(D��o�U��1`?�3?���_gg��7����b�=�٨���n���Ç��g�j���଍f�ք��M�*��@"<wfY�s$s��
g"h�(L"'�,��e��L������{��z :�{�ɐ�ŭA����+�y�,�B���;&����78��3�3�3,�1(k}}�=����'�dW/_�>$Sd>P����,�]w��~����[+��]V��OѶ�_�*�Jl/Lq�5(E���2剚��q�o����@[>=�`�H��"%��r�hr'?��I3`�/.GW	3�Ti�o���&�K�	��?��|��ϱL:j�R�q�0���7"#�J�P		7���RJrU�vdv?��x
	O 
�d$ʘ$T����S�{�����G�s����E����@�o{����+w�cS&�5�|��|!tW��3���}ϣ��G����H\���I���Q�H&�s
w[N���,s2q9�| !���O�h��~������&�E��>�U��& �~^�A�Tر����#���0��(`���������������xc�y
�9���0x�O�͎9®�+|�\fαt)r�:�gQrQ(��90.��ҟ\_7�~t�&S��]sB�+�orb�L�M4x�s2/�>K޽�,y�|eW{�K��b��%V��F��Y��c��	�.H���s�MH��p~N��v����'P���9	&VD`{4�II�l~���'Ă"������4@'N�E� �dz�-//����P��ϑ!Q�;ؽo����{EI= �ZP��W�0K�s~p��h-��͋�P�0  �k� ��)�@�*�4�Z���q�ҋ��a����:FU�6H�%���..s5}�#���/ذ�W��&0:������ڵ1����|%�I��@�_��nf|��0Ĝ�)�݃~Q{g_��@c���@�Mp~�H(B����������.��x3!!a[�l�6R:N�2_���>�W�^e��4�{#�Ͱ�(����p��� -�k��V���d�Ah72d@Lt8`<r�Tf��
Kg�t�GH��$_�<����o�0�Zb�Z�Df��s`9R==zg@_�	10\� C�KI	�S��#��t���.9�ȹk+�����L�-^hrK�^�~�{��D��T��Y�k=h<�[	��ښs�J�q���2j2O��Iy[D�IH8�P^n�[��m��w���J al���	i�>�572��d\8!- �./-i�0����
v|�%$�!��g�Ek&XA"T���8I��D���kN�1�8��WF�,�|@��]raM I��ә�va8B��b��Ť������E��e#�I��|0���l��� �Џ��"S���^D�h�'�>.CeG�s[�4IqJT���\"p=�M�5�Q0��Q�kIHh�Ш.`v���O���td�Ɗ��r��lI`{2W'I��2��m��'�=pޓm�w��S�O�|xa;J�8��ta�0�J�		{ ��0�Y6��.G�����~
Ϛ\����u����1P�P0��AL���";r�fJ-C4����w �s1:Y/b����{��j�ma�c�t��F�}>���@���4�?�f�84*��>���iIt �UN+�f�f�6�p�����������=8c��C ��2�x�\���d2�{}�Isy�8�_�t� ��B�y�Q�cli`�����op{���te�y���7����V(���X�ڹ�}�?wӳ��ʰڎ9���U�a:���N|�+W���ׯ;���7���Hp-t�x��� �v�Vm�\.�º�$b,� B�dr���p��g�g�j(��	9K�-���4����Y��,���y�(�F�R$���<�.(":�$9m'��� J�l�����6�Hxq��3�GGz����%��z$��g02[�M�0a�͏���L�/e��D�L�1�"=�|S42�"�����"�NL	0x=�׀��);%��1,�!��¥�7|VVV؉'P����^}�UdJH�ׂV$ր�u��r�`�Y*�Xb0(T��톛�Ĕ$$$T�ں',MDt��	�������躠<�^�� 1��|��;��W{��� ����/�ka�`� *�r�b�4*/�(�=W��5�U��P�K�yI2������i�b�<:�m��X"���~�����7�b�����}/���{����م��9�k�=��Hd�DVK;iE���s�M6`2��pO��>����w��� {�m��Ǐ�oh@���7�����ɞz�)<��w��%S�sF��������EǱ���;:a�����L.��Y}m<ԕi9!!�f�)�F'ݖ��d`'?�l�?ѯ�������|�#1l5 >�6A���d�D����%F�4�7�O]��6f[%k����ٙ`�*?�wC��vo|���m��&N��p�����'���m�bi�I0�:�)�k!Kͅy܂��魠��G����}�����@{48 �/^D����c?��?�~�a�'��eҋ/�Ȟ}�Y��o|�=��38n!�1(
�c��UخC'b����C�YU�Q u�[��ؚ��9s���O�$��G?��?4\�{=�Ï�?��?c���'����oh���þ�۬�7xv?�j�^���".l�@ot?Az�6�ODX�^D[\�c���B�yo���Tҳ��hv ;8hQ��pgJL��p3aR�(y�e9�9:L�ۈE��$��:I�AQ�y��߃��C鮈��^n�y�(���|\����p������sݣ���'�la1g����󡦟�$ݿ�1�̀�Q����̎Ȕ��Wc�d�ST+жPTRx4�´�]~�[Y�>���M�bQ�klB&^�6a�|�W���ż<�bK�Ƅ�aǏ�d+�G���
�Ŕ��h7,Fz,�6d
�ȺY��[��5�zL��Ƀ�쎨�9m�"}q����V���/���/��WA���sgS�S�/�a|�>j,�@� !?{饗�C=�~�~�}�pL�{����w�����1i�����}�kh���k�a�h��̺�]�a�����,fn�ր��7M�S���o��o�Gy��:u���!'��ϯ�ʯ�9֧?�id`����>�8�����#����f�3#���֔�<���E�i@�A���S��B�QBBB��P;���`�k��[���0ٻm�0�4=�A|r��O��%vhu��^a�b��+�X=w��|%CL?��d�����MNNv����;�[H�����eM�
CT��d��@�},L݅�x���Ɖ\��gv`�B
�B�E���`�:As4s�NMS�<q�B1i;Kf�_ZZd�®?�	��z�bR��q�&-�ǥhо�~0��7c.��$Y� i���4��/�"�Ї>�ǧ.w�d�����}�c�+_�
��?�c����_Gf�Ra��l{��qB� �80��1`&��������"�4�fE?��f�G�_��_gO>�$�������r�Ѓ�e_���q�q��\w"�nW�K@(7Pr�JHH� �#e�#!"eT��@��rMӨ��� g^ 𗗗����������KLi��(��!]b$��f�,%�J��7i8����R�_�F��"dњ,�:���t%A4�Z]B�ǌ0j\�����ܘe���)Xi�`���M*���I�Ϙ�p�g��
]v���ٴ�i�ߦ�AE�"M���k��>��#MM
�����t9;}�42,�����`��q��4i?n;�JZPـs�G>�l<EÂ�ΣD8���HF���ym	ا�6hp|?D.����HI�n3��Ѭ�h8R������ј8؄�����IRl4 SM�-�yFZ^��L���������vZ���B_or���Ѝ�b!�.0;p4 @hCD`v�P�7Q����;,��#vz�v���&U6H���)�9	��x�3N��ۚN����U&������mj�o]ӁH2e9�����~��я#�)Äe�?{o�+I�Uo7w��L��Y�U]CW7���>���"o ��H������ 		$��@b��j议��̪�3��|0�l�m�a�'Δ�l�"O��>�e{�����  e��^#�ت!�_D$�q��'5-u�\����tlnn����V����<S x�]"[�O/��A�7�1����� �����ү�گ�8<�y�KOO@P�A� ��a�n��/�"���P�ƀ����׵�Q�q�y��������y�ba�l|�G{�E˗<CI�v��Y�Hx�_G�	��Z���>�TŸ�aΐA1���� �J���iP��֗��3��-G%Df��\�pܪ���E�2��Ia���E/}r�% �� 	�'Xܕ�I���x�J����Ѥ���y@����_��_�k���P|��c"jN��r���K-E K�f����0��M��t��:<:t
\9�` ��Fk���9qU_�}��ZVM+U7o��h#�6�E>�|/���֭ۼ|����.=��jww��B&� �z=�yoH�	���T��gS���n�c�[Է�KM?��=~Dۏ�� ���qC ���I��?����0_�����mz���a�˫1��qӧ)�c���En,T���W���]���p��*J�j���W�E ���.?�+��+�c?�c�MO�Xr�M�C1�W<~�'�~��~�~�7~�Y��yb?F��=B*���\�}O@��	� �@�T0:�/(�c��T 0�P<�i���,�y������_�ׯvB#F��z�s|*��;O���d�`��!IE�����������m�A��?��+p�9�וK�{<c���I�����kt��ν@�޵ ��}�s�ڄ��0��ڒ��P�B��CY����)k%� $�H~�t�|����__� �� �ͫ��b+׎�V����X�v;�no�󎽽M�nQ9+��o���{l���9ծ4�킲U�u,�嬓/���. a�Y��L�}j!Tt.��۰|��U�`ճKҝ�'��f�cl� D�P�xUY�K�)�����m3�
���h<�,_U@�ڧ ��+#ܒt
 h��Q�����	�F�7O��Uh��*F��+_s�-1bĈqy#��s����YP�E�6>��k7�X�:��=�EG��ľ>9�LyM�����k�AK��Xp=j��,���\�s0����?��������k_۵�beߋ��BT
[�]).�NW���Ƒ;UŌ����W@�5|���NNv0�<^�Xp���U���<���T��3jeoh!sjY5�b>���u��0?�^Z	o�%�?��$0���گZ&����M_�+�>h�
�� 2�}1���{�~�g����o1=�\�
m�_t�xj �
Ȗd��o����Lؓ���J�i,����O������^*�.��9�79�G0�W#Vi�'��#Ƶ�P�-E�3���-�K���+9 ˊG�ao��Tu%�҃>Q�2����j*íS����	_)y/����	�p4d�ZTC��)�z�d,��O���֯������D�6D�e�r
�-����Loߩ�X�D� �s��;���#����6����s��д*,�l~E��]FN��#�
�]�5�cx��6G8 ��y{��@��c�1�;=�.i�ީ�k�H퐒fB:ƫ3`�-�.��=���3%����s�_��H�i�� ������ �D���aw���oHe�r�~���j���˷���\4�I�_���J>���}�"����u<�����`������ �@Q� ��ɍvfj@�ؑS!@i�Rr�/x<� '1άǸ�-��4�<.�e4���Y��9E��􄺙#-��(�3-�/�N'ňqM�;T�Ӂr$+*�؟G��y|�s��y}�����uM7�%����$�q���P�\啱�y��' �:u2��>�y�&��Z+�i�~f̟���r��oM(����t�&��K@Z� !�Q��쬲����.�5Q���SK�� q��h8ත�h�Ռ�(y\�ݝ����&�P�B���`m�-W��ۿ�4a ���FY�h�7����-@f=n�ºCrX�r��{�.ݳ����:��3샛[�;�՜�[���$4Z�P9�36���s�eج�>W��q����y|�k��bNNx�2\j�Jf�%ؤq:�ίM�1���������e�&i�v�|x��Ϸ�_����;|<'�)���ޝne�s��=��6����U�دO���.�Ĉޯ$�< �h������A�}oz���B��U$�������(�zЮ/�-���˧�#�r��u[�0V�bĸ�����|[�ku��Ｑ������u*��Jt�Mk� �۱���Rfo&)'s&�&��^��P[��R�H��TX ��<hcs�^�s�6�6y�GG���`ς��#��[�����C��Ex�����[ 	��3�Ă�n/��������^$�Hd�� ���]��L����7^���	>ڞT��&��s�V|���-V+�3�X��	�m�&(�gz�֓�<��G\9� yj��� ��� 0K�w`�P]��HS�yq�E;�2(i����w����Y���n#�A�Rts:/�$T5 *P� �A���<��� p�R* ��`����b�����Ί6H��(
�!���F8���#��pv%r@bĈq������,r�C�t�
O  �r�\��iB����῁��[i���F�Y�p�;�g��$�
E�3�����ݺsW�Szà�0 �yU�n˘xn��ӭ�[L�*���+ �AF�[�$��:��F��etk��6F���Fo��tr��@ذB{*Ai�h�Э�2�)O^kn�R\��%Ts�}	#=��)N��v������Z��+K��1�� H��-N���}���2���yC�n��N �X>��i�D|�� �S�|��̀���a���Kz���K�bá
��ym�s˛~��@��M1b\�Ё�z�1b\�`�� ��&$ŝ��T@t�r��Ms������:߇�L&JOh������O���U �ۿ6/J53�-��C ���el�.FȲ _�4�Θ>];�C�VI��njQ��*�PYWM�O,���@b�L,��4�~��&���ŀ ���6�m@���(%K7�J
fѡ�Pbsǒs��ۯ�蠭7�/�[�����\��W�m���$�7��:�>w=�TĐ�C�yUμ�-����<�_�7��3�������FZ���	@<�"d��+��?.n�X@��ۦ�Ή��#-m�W:T���~����rk6���h���������H��$D�0�7���0�����ԬV��@o<俗��N��&��A�K�L�L�w�
A�20SV̼O��u׺�{�Y7]�����1b�xv���*l�h�sHI�<�l���؁p̗��ˤJ���ę���F>ޛЬ�s�3����p@��M�SicI{�+���HH�*a�n*���vs�9�4�;uGC�j�N�n�>/$oV�bW�������3��3�����uQ1o}�	_~�^N�_plS�L�t� _cb���ŷ��<_�I�tYQn��J�~�=��Sb�sjf�|�JL�~�N<�^��	�L�Ʉ&����9�X���غ%�߂�a����$�cb�A �� �ԊE˓��ƾ��= g�S~��s�O��b򟥣��! �ѷ>��L|� L�I����q��' t�XH^�� 0(:O_X�R���
�������y�˺������A_fx�;N���'d&�]� F���@�g��ǈ#�e������5�瘡G�gpTЖ�����S��� $�����ٜ�& �@l���Lp@��ר_��g���p-�	$�6Wb�_�{1�B��$R<���$��v��bW$� (L��y���_�,��T@��%.�I�rYD�~ֳ��(�H�
]�sw��6U����U%�#q�m�ImU)�K2מ�e�ʄ��TM8w�mc b��`��"(t�����o��oY��Jȩ��(pB���F��@��}�^����
X�����O@N|9*@C�T|��'�5,��u�e�A��?�#��?�s�/��}@<��W_^v`��Ag*9)<I���7%��w�^#F��5�0�c"w $7%�`�H�M ���N���T���gB�Ҕߏ�3��[����k����,Z�8���<:Sb�ke�E�0�¤��Ԥ�t�Cb�I�)(G���N��0���v.�-����;;�:��0p+O�rP} �e^�i:s%��0��i�M@kV���-昔�n���4�E�6���x8K{�}c�ʹ�[7�~���0S�߈�
rf�;�'B?��?J?�?�d xVx(���g��_��[��N��`�/*�L $р� �����_��_��"��`TuJQ;:�����������7�h���)}����0y1�V7��,��]��>���1b��P'܏#Ƌ���]�$HI�VL�9�O�-�u��6�<&�{MB��a�w�ث$1�$,\��d)��w'��e6	Ǽ<ZTaH�\���H짍WGQ�i<��H���z*w@�n�'h�
�bE*�Y�
�Ĺ��̣���vy*��XP�Ki3�T@���%ǸV/����w�x�)�m]]b ĥ����X�(�"�M1��4�kǧJ�-e~Jk���Q,}���_W�6�D�M�]�H�9a����V�xoNŷ�e2���&�[�3-|��������.���&�v����؏ B Z������7�M�h�:o<5 �_gD���Ͱ�?��?�H��8-8x̬y�,"�2�����>��o�6���{\.�ʃ��;|{}���jP����>#$��o� hͲq��:̤��D9yg���A!N�L��b\���esZm+qi=T�9�z_�օ�9i�R�N"u����#�M�ԅ�P����0[̍;�8QC�)Op5�f��R�-Wf�u�.s��|�&��������UnS�IgΧ-E���
*R2��D����v�Po}}��ݽG�рf $��
&M"���6&f�%P�R4�����
V�2��� ��Y)��)���ims��#C�iϹCg����E���d�dq!�j\;X�ن�i-��\��6 p5І?�L���>��a�~�*�6��f�����`*a� �cٹ]�®hU�TM���4�s��Ufi�snm^H�'A���I0��Ha����F�W�h�t,e~I���w.˻���U���ys��%Ucd�AND�D�^mxڽ���'9����y���������~�W�sk���fc��6A����ϿL��O��=z��A��Cy5�����m%Byj ��pv���CihU�w�y���p(�
�"�Ob�}l���������_��_3c��ᓔy�<T�T�{=χ������������ӏ��
G�#�5������xh�"����_��S������k6�9�7��~R�� �Rz�u��C��GEI7*  �'nB�I(?M'��������[[4�w�ud��O�r�e���À	�Ll�$�ͷ�@�6�fb7�G9p!��PO�2�HJ�@��� P�2��z�J�� �0��2�vv�����x�&�cnA[�hs}@����h��Tz�i{{����oܲ�I����,�)�SL���>ۿS�YpS�j(~a0��T��U%��kUs�����T����V��RI�,c�лfyo�yܢbxY&Ҽ���!��o���t��=Z[[��\���K� �F^�������GpB ��?���]�:rR� �LZ�˝wܯ��R_���P`�_{�5���z���
Yh���7�I�WE��{�ǟ��=�>����Яz���	1b�$Y>V�d���5�#F��a��u����'�����S%2;�tF��?����.���]ι%����t�ǁĽ���������e)���;�ܥ��!=����Gߢ#���C��(teL�wh��O�h�Wκ@F����Zs�HFQ�@^������m} �����]n�?���JFF5��uZ϶����:�9L�鰞�����紷H���{�������ʎ�l<g?���n3�ٛ]O����]�d,Fy ��f<�6�j��o ��*��+D�N6�K��J�YỆ �������M��W�B��˿L?�c?�]K�v>��>5ڿ����>>�W�mZ�����s���n�wX��
�~|�#_@J���������Ƹ�� �B�������a���/6��hWAB�qe cĸ*�g8Ë�:�T���cĈq�"�~�3銮�G�v�t̴�O�bP����PU�$�uI{���t:n=��=1�K��g�`�v���;w�g�t>�r���]��i�|K��r80�״m����'���I&������ji"ٷ� 0���L�H�-Xڙ*'��m�0�^����6�)�:f��KhkС>��'��t�i���̮{GU����-W�$��b�}/C��N3�
�㪓��X�W� �]~E󢤉��\ ��ۀ��`�ƍ�=����d�&��O�Ҿ�
�+� �?��?c�K��K�S?�S̵���OA� ��p���_����w�L�+�+iہsR��vX�_�A��)��O��O������K?��?�+�-p<�7�-W�)�}��=�8/��ĝqy�r�1�F��H�.x)��Yͳ�b��i2�>��ŸJ!�]�T,� #䁤-����@$F����҂��x]q��~缶�J�B�+�~R3���gؠK�Q����'��=~�M���oҠס/��6�7�F�l��m�ǹ�y��o�z�6u��o��Z �O�iI_��m�=�-��2q9��<��U��@��`���V��:��I����~�[j�����|εmg:��
V�|ER���9+��,^�1g��k�l��ڈ���=�X��]�����.4;�W%Z����4�[p13ª2L��C�ǷM�����[_��������p~D��MƳ�%Ɗs:4u��iM�]���%���#�F>r4@{�}��[�E����O_�җx�P%�X��ۿ�w$���Ϣ]������ Nʳ�f�W7l? 	۠<�œ`����l( ��|���������ꈗ~[���گb�%F�1b�8;t�{�	��]�J��%�E�* S2J6��%���[��?, A�90�<Ԫ0K-*Y�&�J��!W�-  ��T�Aϩ�_��(x$ j;�9*/ 刺�r��<��pmg'� �ɂI������v���$�uQ2��F�7pD�bʊ^��>O��L�v�ŉ#��q��F�c38+�F&�\���B�`���d�3�xޤ9��z��n߱�%��u�I0<��b���5_,�o����
��{~ Б����"�S9f�8�O]A�_	�������slR0��l,7TA¶.? ��l��C��.�B1b�p�8f�B���ƈ�f�*�q]Z\�� ��
F|�eL�t������~�������z��q�ڧnV�O��EU�cy��.Y�2X��+��5B9��CT<�Ѕ�Aa
��  P5�a�@]�
m{nUQE�� ��p��ݕ�ǘXF+�g��f6�� V� F� ���$��p��d]=O��N�P����,�8Y`�
8+��e�]gP�1��� �<��=|�O?L�A�:y��:�R
H�Qu���� ��� t���W�3H���ȳ�z&N�O\�!d�c�}(�`��#�` ��f�����6�� �ń�%d�R6���U9[!11-�qM�Qщ#ƕ>��k�Kz��>`wl��:��Ua��<�O�/tF	;IY���p�Fo���=����wޢ���9s-��6Ja&��vW��E��&���8����X��k��)�)���0K��%�m t��:�-��p���y�  /E-@�E(�v�F����HH�C�h � z*��pNP��3�u��\�%�(u��N\uE3�3ZL
�o�1��Il�7�&&�w�������i}��@�a"���ZY�a��%���	� ��P��r�Ϸ����`��0�ȻQ��JgU���Dz�w6]0:��& �+gBM��h� �����a�{�vv�2��'��~`�mI @���h��y�'�gc�B��6{4{��r�wv6'��7v�V�/F����b?{Zx ��	��Bw/���[j'�Y0v�%{b35ň��>I*3ђ@\$⋑����f����#)���/�&��$S��&���7->c.G�;���~{k��Ҷ�V�,��pp��n�Ni�F�ۡR�1@ ���$"��d_�Y��rI�D�6��Kȕ�2$�,9[���<k�(T�w���]�u�0�k�;�
�����}�08��i՜U�jE�u� ~?��{���C�S��d�]$����r�RBx�$KD�V
�^Ǝ�����\k��)Ԝ����Q�ߧ}�us;F��j�^
�=Z�@�<U3�'��/_WW��i��Ů��k��T#�9�7rl?���{���!���w�_>|�$�i^�+a��r�B��b��{7s�'[1yș���@�
���M�u\��rlF�.�-�h>9���1�n�fzܱrl)%tǈq�B��\�ۮ璼�y�8��WΈ0oP��E���sE���������X�C�M��є��>e��%��Ծ^;��:���#$����,���������$�kL�4���?bP(�1Y7I��^��B;�1���$����ى�c,UH���D�|��ϧ����S���m����<6�����X��{<_�
mV6�LRQԪ��f� }��]�~o�|ڞ0����@���θ�V
X�y�W�
�w5=E>���U<��*?�����=��VX���q�6�������e1bĸ��=��*�¤�낎�{���Mif��LeϏ��h2P@r �7f��ȍ�$  �Z��	��^��v�(I1������]qo'˫Q�49\`�h85K�u������0���>�D��"�9ڞ�SF�f5/�i�D)+�d�:�3<6�C%IeF	�!�Dʊ�r�	�����ͻ ������.�א���b.gi�����s��\(�n��^'�+��K@`>�G��eYӃvQ�']ϧ]���U�qx�1nj���	����)St�L��h��Lڲ@�P�	�:�.������E��4U�"�
P��S����*���	WER�E`�j�Z��sp�bz���,��mN�U����J�T.pʦ��	���d1�ץw9_c>�+e�z��M�j�b<�~	��l���VKci) P)*��[���d��7�*F�X�*�A�� l�h��L5�����i���Uҹ!��!0�O�v���O��Pi˯z+Y������
�g�+A��ď���� ��H��u�G�p��-���M��_�ܧ1.G� 	Cd�k��%�u3�i-ki���c�s�b0wBH�/��eB���O�88�Yj~�3P�,~
�1�O�:P-���8T22��I��8���y?�"���j
�Z�� ������� ��L�} )��c��ؤЂ$�V����!��{�4ᇘ���$mޮ�O6�*�Æ����N%
a�[[�h���J��:%0a�e�━SQy��|����˪��-T��!�:���C��P�B���<��{<oÏI�r�������.'oh)큫��g^�
�\��cĈ#F�7/$i^~���|�J�1��WT�M�� |�ß�w{�8�=G,Y+�U�3��OH�"e�*�R��$	P�����<��E򏲆�f˴؄0��N�>�W�ӥ5^z��K�����P|��d��� ����/Q��;�_�۲����	/�Z�؉�R'A�Z@�&F���'n$ 9+.��H�W%���F%';a����+F��:@��r�cN])�̩�ʥΠ�4ͳ���n	��$�uQ8�G�d�x-�U� /W��	�܋����PP�������.�*[��U�D �>A2�8@���}��2(I��9��q���)��C�M�=i:b���k�Ը_q[2b}8�nt��w�^�I��┼ �����~x�� mۋ���~���+/��j��$8�c>��D�7���	&(�;��iQ_�q*F�K&Y�VF�N���/�"*b].!6�Ź̜���
$uY�:�*gs�Q�S�$pDj�A����^���9�,E�jN�X�,�@[w[m���ܧ����B
�	�(��.� êP�YH��7i��7�9�V�d9���|ZžT/W@����˓V�5�y/���O���
� -��O��d��
�Sd&�k�=+�*�e��<�x��g=�e��i��L~��Ίn�@5�b(�
_���,���U�\Ly��Ah_�1!��죡�%�g�U�2q��bx��~r�o4"��i��s��#�E«4�A�v��mxf]�Ԯ��|],��WD/��ȏ����/��K&�n����I�ޝ�9��@�	V�`��yzho#^ޠף�ф*W�Hs|8)cV�Jx(� x��JS!yE�P�I���,�+�$����oY��/�J�^	;���]V�qU u`�w�h�������i8ym� ��ƹt��'˓_\ut�Y(-�$��v�ƏwۇDZ�*#f^����Nָ��2��=� �P���Qp�"���i��׻�7�W�������p�y-}枛!g����?I�U�6(��2�����ȟWú� ~�{$�q�����Q'��/:�;�l3?1b�~�>��y�'wƈ�EhȞN=i% %a}���VtY��O23���r��b2C�oo�ҵ%��!d�Ĭ�>Od�Y��V���� �@eÏ?F6C�$�n��*q,���d��S	D1 �Ƌ>)��+�BiִY���>�/�Yݼg�J�Lz6A�䦑�^��pR1�ST�����̭���`Ϸا���s�SF������\���V@"�x����1�phw��ѻ�FOɱ�Y2Y�蟷"H�1b����?f�k-��uY�j���Q����)T�����=e�wgd��L�w���/�Ym��r%�T�a���MeGD������h_�X� �K �ܺ�2<	{͵XU�D��s ߕ5�'�:x�Dʗ?V���B�	c�
�xlǿ�)�%̽�1�z�q^'��!�� ���D8k����Qy$F��-�B˜i��?!Bwhw�&�)��s�J 9��'eX֜����Ƿq��ˠe��暸��[�PM�.�'��w�-�\���d��㷯�����|������LDo;��ĸuJ*4a�`���89��{[�]��d{!��,ϸ�ĭd�|�u�x�t�e�S�{}_X�{�6.�~ca���/^[x����$�2Q�0��-|@(0̡1�O$�)�,'��8r�UK�(�eň��C7���9d��~%�\9u��'�^W.��+dgozx0R�p0�v������LZ�j���d�5=�/H/��9��RS���r[��]}�ddS'�++Ya��s�!�H�/)^��y��lD�ڭ�R�k��D�"QÈoy��+ߞO��}xRy� ��=�
H���q|�7�C�81"��P��S1��p>���������Xp%ˍ	���*d��D^�-�)�㓼yB�� �%�X���{�bĈ��+�,U��1�vh'$�Imr2�0Q@����HCb\'���C� 9g0I\w^,��t�)�)� ��d�n�����eIlh�罦�PW�%�θ/M��]��[Ujj��Fk�Q�|]�	9��v�n�W�ޘ��Lg�܂�T[v����N&�t�L��BϦ�0 �ãCv��N&�z#;n}$5 �D���Ą/,^�
�u�%՟�E|跴�cĸ�J0��1bĸ�����9r3�i�%&V@��}�*	�r�2��r�Gr�p8�x�+�ƄD�bH�!���jT�Ԣ���8�:�u�t#��ElZW��*���@!(2�	��NʫO	bI�%�u��I{ �O: n<����c���/�s%�Wf�:W��%m�_I������2��j���}�Jn_�N��������hb��p�A_���<�p�s'dd�D �*Ċ��U�5�B����UL�T�1b<�X�ԥ����{�C�E�]�z�������g���j���p���: ��y�O�@2v:��|^R�31��C�$�PblS�h����D��e����[�2,)�WDR,( z�:]'������,כ%�nj�ț4 D�f��Ʋ��FVƘ����q-�ȃc��&.�)�$���
��J�Nठ�
�������PyR���08x���Y��`����ʖ�&���ç�B� ���q��b�����hKvn��X�|��8���G�|?�d^s��>�L���]�v�70']�uܥ��C��ۿ�>)�}|1b	��J�rƈq}bA��Ap
���&�";��������/��R�0'�Ү�8�;J.k��HZ������k�$wRV^*�3����۱DB�۷_c^�h������:��t2w�	�#�����}�^sqR!���(Vl�N�6��� 8(����<�>��K�\�a����a�^�1D�g��ur"W��A�MR���uYT"��� ��L@�Z���)�&S:���|lsc��6����[��NA�fv��]��ߓB�B�GZ��j@�����]��1/#���s:������x�`��꤫�N�W-��>+�T1b�x��T@O�	а׫�&�.t���-�Aտ�,�Zs�����Mӊ�2�$�HM�G��hx����w�h�?�,�A�zn�Y�����H A�M�AJw�K�>+*�u+A,����KCa{x]�y��a����2����
[�@��,B�N��@�'x7�`�߈bI���n�<Y~���o~󛴿'�c��w
�ϓ�QI��b�M%�\�a�AsK*��a㸏'N�]��b��U@b\,��b�)7�{�uXӎ��y*�W��#�u$m��BtT�̈G1�s\Ǒ��z�}���i���.}���t��m��KN����U����6�f]6��<��r�Ѣ+K�v�2��]�H��*4�ڗ�ޟ$�ƀ0�c�^-��ҲYr�M��Cy�T����X,��H����r���'�g���X��p� ��L��_�Ek�k����2ٟh��y���ļ���Y $i��q�8�D���Ƹ���؀�c�(Ĉq9Bf��߳��&�2����0A>��x	�O(4}�;��������666(���Ν;4�x�܆���h#�Π2�Z�P��/����x�C]/W@����v��7%�Q����q te.� \)s��ک�-��5�T��qJ�-\ރ�o�:���>����w�h|�65��d<��Oo����;�R����i8Q���<��4�����BҊ8u��Λxҏ�q_���#�z-��,Nℬ�89�9���>3K̩�\��;yY�k�E9:�nc\��=�~fkU��T.�;�B��1#F��P"�ꊏKp�>#*"Yޣ��H��t��}~[x��QP������������ï�?��8ͻ���NkkC;���P���$��v�r�ک@��la �   �[��ù���,\�ܮ��A�1��������j��]�9 - �Mk) гC�[^ں���bL�>¡���������4UU�>���������c���9T��v{�v]s��Y�`�/�{÷�.l�ި�'O�Z�c�������hp�[U�����
��x�&W�p��cE��Y�ڷ`Q 1�fx����Y&�q7�� ��X���DhZ���)��\AR^�8lq���`L����AB%�w�vx'�$9�Yx�x��8���qI�dM�gCSA �r�~m~��'a�D�ʚ�LT����C8R��_�c�L0�k��M�䰑����D��[�_U"v��`��J,�:a{c<����8��d�V�s#���*��m���8@N[.�trz,�7yE�b\�0��L-P^`�(�#ƕ����#E�8=�3ǣ��P������"Ř~�����J&�ռ��9s����Z�Ԛg�ۓ�IsD�>��sKXY.f�U��x�V�/��`�
�����Vɲ˄�Ti��b�畗��m���?�J%�]Yj�B��x<��x����ë��1��*L� �9<ඬ����L�2q~�q& q�9B�cq��iI�='˚�K'VɊ3J1�b��FB�<�13]�ܧS��cĈ��c�Z�]̈́'�I� �ݶϐ-m�������6��F6ٿC���l�7��kk�y��7�{���ۛ�~�Z��G3ʲ'�hgA;��9�����wrr�:ϐ��ˀ÷H�-K�9�MT��U��-Sh �X,0�6�^L&K��{�Mz�fx>WcR����e��a��S�|�7|N��2 ������>�����{�����҂�Ҕ����� ��JqK��g��|���G	-�ޥ��y�������=n���}=����8?�	@쎚`��;�M�e$�/-�4_%�4�
y��j��C��K�Z��'�S�ʢ�A���9@�Tu7|O0�}<��b��0���-w'w�*;��떡nƹ&F��h���:Gp����溶8rc�9�]��!,�k��/\M�	�Z���&\�k�o#�uɺ�2�EI��nݾC�N�&�b�sݠK[��я���C��������G�%||=�)��j�0\^���?�`&�3I�[-P���l���7Qٲ,nf3GCK.�Is6GDx������2� 9<�~�}�p�.�M��uVyS��:��#mU}���N�A�~�)=�~��V?�޽�
X �{�����5H���n�^5��@�Ա�4q�e�&��B� �0�t�i�����"��aK�|�����Y=�~	�(�#��*��jT *t��C* M�V�W,X�W>������/���TL�;�bm<F��(�}�N�.5�g��#����ʔ�e�w�CS]d,`Pv��0s��r��LRڼu��������?b�묂5�J��1� @Ա%I܅ ���u+�ow��@��3�V,���L����ȝ��?v_A%'MA ��ZAFH��PW�qX����4��lZ�W��U�F\�	e��Y���m��n{⤄ö`�&1���-��u;eN�E����+ tCȪ~����O��M:�ƸIq��4�����U�1�u,T�㦴��Ea�t�`�O���D�� h��t��u��f}��d5'���'mG�'�5?g��q
� %,h�n��[���o��tp(Wɒ���(}<]-��Y���z�t�H��.�����U������/�f8:��
Ե��HQ���a�+���ubo��5��bpM�ȍ�"̅��y�ĸ��{c����	�B��ňq�#] �En�J�2� e',�ĳ�~Ͼ����#��ާ�M�1k��Fe�����F��a$���lb��,�͏�a$4&D���s���oQK-X����v������'�9�ARS�r)o��
L͠J ��h�U��� 19�hBE�(P���}n(�ˍSH���������Ą����"�l��Bl�ӗI9�{�\$c���9i@W�ete�c�85��6RDW��^�ܩ�$7��#ƥVZʒ�����k����mBw��r���l�A�k׺>�cYL� DC�dńmW�P�j� @�Ih�*�m^�4���֙^��vU;�(%�DB	Z�¨Vp Nn�3���L��� �%x�N|�B�?.�{��eOX<�.�'������hqͨ-��C�ʂ�9Zݎyp$�	�ƄpeB�-i[3���Y
��+)sd��Y&�_L�0�Q�T���=��r<�hyB�Z�/�1b\���|�L� Њ�9>�Ǫ_��:�|�꥿Vs�!׳EQ�)@���Ir�4�iA	�&��$�:�	J�\�k����r+>G���Ӂ�Y	�n&���B4c�cI����׍>�v��-Q��u�mH4�e��01_<@B!C���Gl�:%^����H_�q�C�n��YVK'�h^#�͊���R�j�u�����U�Q�\T7� D�RfkV�\	Y�]�T�v�~u�e�,�r�"Q�c1�a"� B�6*�	� f߳�������K�n/�	�Tq��ǪQX��1����jYyׂ����D([�'�^r����{#�W0�zV;g��c�8:z~ĈqY#9���'�o�B\;��$�)����Pg�yr���؃��p��~5���(\Ѯ�"�+�[O�����*f��g'��]�89N�T+�isBڕ��벬J��=��W�d	��v�}"0.LӼ�>�V�#L�эvm�.N .g�O�_��'9����}m��js#��j���T�k�u ���W�R��H�#�#��S{���!���5�M�Ħ��K�t���1b���u=���1oI�MPȻΝ�.)�{�*�y;}h�g���P�>�Ț��#W0xC�W���JT�:��
��s�(w;��)��7\)�]3�Iricmr��Sy���g= ����YJ�ۂ ���B<xL����^n҂,p�9�,%���|�Õp�ZY~�/?Β��6�2�_a� �^�J���5L�g���{}�<�P��:M�N�'�c?�؃;1��,g���U����/I7U$'�K��Ir�0{l�Z]f�=�r�U9�?VW~�'�/��^����D�ӄQB
S����ls;��QN� $�u�X��9����Y�U�<?cd��ݷ�iW �v}���7m�}jXE! ���So0�dx��$zH��6�6y�	j�r%�M5��E�|��0�]/L"��K�)Gz����e��eV�S���U��S�H 'nى(�z9AM�1��z$���dRȺBF�F��]�n츂Sn�x<�έA��l�7"��f��nn9Wu��Ҷ��x������y�������Mh?<OD ��MLR��p�A9 1�G����#F��^m�*+�q<�f�X�ϰ������tB}����+4����O\�=|D�(�@Rp�-[����s)�������n��7b��,Wo���u�z��$�t_��ji K��f�����9(- 0�X��~#v!��	ݾs���n�t:e ��>M��V�٘>�η������G#^7H�/�����ڼ� �c�3v4�v�/>Λ1ǟ�`Y��$p�p=�(m��Gq�8����#�Տ��#�,[Kk
nh1Ml%&(b- �ze�F�4����}���i��+# *� ���@P��~��PZ��j\�!���_�w���|]���O����D?��������;�f}�����n�>M��c��5I{8>r Dںnm��ud�F��������e�1���c2���!M&���m~~����DQtxxH4׹8�s�ILi/C��AX�]����,�e�ݔ~U�Lg[�e��L>� ��Meѽ�4d|�	vb�x��Z��+��'�g���ҽj]�"܎�r�����~$��dK�s��&��keY��r� ]-�}�6�]�0؄y�3���&�[��$Y����k_�����ttx�gI���DU���$��%kkkt���u�����f3z��}��g\q/B�*���
��U��t�a�#�c]Ъ䕻�ۇ�' ��������/�_��O?�O�x����O���Wn�l �CX��l��n�~���{���޽k�؀��������G�m��(X ��������Wn�pch�5���5`͏nw_y���&������������ �0/}��섖�,b�%�/�P#Ƶ��P*rCbĸz��e�rf@|����Hp3̴�$�ij��>�:��ԙ�(�c�II��#�`o���mo�X�Q3`��ϣ�O�Y[_�w�~�^}�U~������C@��3�H�Ӂ� 0 	  ����V��,�j�OL};�J��D�|��$�� Z��l�������Gt����Иb9@0 `cK8��tgg�����/x[o?���G�m����Y��t%�յ'��_
**���qa��F4V�^l<1 Ib��L�Ձ5�1�R�V�
�����̗,�#F��HиE���$U}H�#&r߆�mk�/��u��vy&����k>J�����4Pd�(�p(��C)
�D�tB�M�<��lJG�6�ߥ
�S�Iś����<-�"�׊&����D��ɉ��^&ʭnA��)b��bFe9g@�	�a����e4�T�*#w�nY@��11��T��S����x����s�`k��j�;+��H��'� ����*X�c��~��GߡH��"BD�1nJ���fNcĈq���EآՀ�P���F1H�����& �]:�zr~�K�Q���k*�)��g4�`!GROZ�
�4l2=\�tvD�nNs�>�̔M�S;�<d�`���n��F�-���C���Q�9u{)e%H�<�	�]^&w$���C�ပ��Z���Ǐ�t:��G���/N]x*x�ה�ѐ�v���ޤ^?��)�M�-;�M�j^�+�|�ul�>��b�M��z�{��q���*B����n����ƀ[����r�n�`g�[1�uD��Uze�ȓ�O"ٟ��'A�_<�����{��88A [
>y}5�ɤ'�mTu]������ּ���)�eA&O��X���C�/��YʁYYӞ�w�%,��X>q��+�(�H�xLĈ�r�{X�8J���db��ڪ| ��"\JH�&)_��ׁ{ojgD���uӟ�.����b]}
���heV�x|��~Po��e��F" ��yE9���}z���SM]��P=;���u!P���]�w�5X R��a��.taK�Rڸ5��l��[���'��|�������eAC��u.�JOm��Z[�4�3�0J��hy��766�o� �Z�ݞ]CU1�4����}e�:v�zy/h��:���7�d 2X�<ZͲ�0�*>ꢲ�i}kdAEB룞oS���wib�m2��1��=��#z�>��@�s�%gլ:���8R�|��o�9�%���ҙ��%���D��y�y&�j���\� 謪��j��X95�ɓg?�;C��fq��7XYL������-�6�c�18��|��>�� ��u����b9'��\�Pf��`����6��h������m��M*7ێ�Gq�ƍRq8��91s/F#��+��6��` ��̣m+��l��0?� �v-O�}@���_�۷7- ��dи�#@T� �{m�F��o~����LX�;wn�e�l������Y��K�+(^M-_��������-pX#���i��h����`�5��:�Ohj�c|d����xeb��J�Z2��L�l�cE�N/��s7���!{}̊�}I �@���IE��5�`�����i�A��N�)g����,/|���KJn8&9�H�x�@y/��ul��q�C/��Y�1-s@�$F��'�K@cт|���ǯ� �c6*XY*|L��g��)����x63��m��x��Q��p���w-��0�TA>R�6�fl��^Ŝ��[��P��M� Z'Q
(B+��`İ_�+ں{�6�6l�Jt;R�r7 %��e>Jm�_1�Ĉ�Wkr�eI`�gm�.+�v-v&`�*Q��[�T��	���=� !�F�if�Ui��j���'L��#��S�ߏꍘVܦU4`a+��6]�0�oR�� ��Q��#<ɚ��򼟽L�@�g�?q���w�=i��+�	J�1�G�#F�K8kwi'E�p�T@TZ7��Ư�q*R�X&���x�洱v��4������<X @��F���Ǩ~@�M�\bm�9\_�$�6 @����Ɠ1�Q5�����<����u1J<Hr�� u��.���W �kت$a� p���Iӎ]f���1i<�J���2� d�B�,��R&��Z�mb��t�|^�lVp%�hG�'��7�}�j����j���,�ct'���c۶m;���ƶm��ضmnl���N����ӯ���33]SߪO��.�A�H=B=�^�[�ɾ�h(�!�0��=d��5 �k�������r�����׺��G��o�F�hPnG���d��?�1��m�e���b��ÁY�wM������R����X���<�z6y�e�AUKku��3\�^���h\�8KWr`�F:�B}]:���^y��.��O=3w-���	����ل��� �:]�$�-2¯�P�����������"�!�3(���5����[��:ܕ5�1,p�M��trCB�f�dO N(^��=�&��9�9n�d<B��CTϜE�溛�|�.B��:\�L��c�{N��ߞ�������dA�{Q`N� �ڰ��*�E�����V�H@S")Z���5���󇶚�����M �%�l�|��}�Ʃ��ƞ����	�����|�y,<�
L�k@w��7��ć1U���qYn�~������;�wvH!���#�4;�'��x�Fd�1sڇ�S��ϓ�&��w�{Ϻ@���3t+Dwc�����d�!������ ZY�I�דh|�C2e~J��+����6`,Ap���d�U�|�<���t��f�lM�@��6
���"y{i�Ԓ�I�Uko�[v�:���/�>���b��km��s^J6�.89{T��vP!Y
�ї��Ơ'�3JW��~'�+�y6ErEs�(��I
8�*w3�V��MD���d�
Q��Җv���/�U[mYO�/2΍�fi-0n��ï5�,�`�G=�O9y8z׵2�%�=b�Z�lZ	m8�S��F%꠻�j�%���=H1r���*x_=�o�윜3��lNW���\�x�ēA��<���^��E�uE�@�܁��&-�mɄ���梧<8�Lv<����J#�b�6JJg��aTB�ժ�d_�FD����L"	G��VNg��X������ch��W@��F���ĀK J�j��;,��1��Z:�7EB���2��Hi��z�vԱ����y!��i�Q>�Q�D�޴�aԪ��qpk��|����I�\����ZCE��|��)g9�?�60s�q6f@��.�$Bfz<|꫉�����T�Y���W�m >s����@�HҊc���{�`
:��������5���z�t��~Ȇ��F��P=17�`T6d���4��vp��2�J%�Z�C�8���A�����na�.+�7ru$�9�Ó��RL�+�~�����7��e���%��=M@o�N��W|	w� Ë_.��nE�C�pNt��9�Hz'�CT8�B�	�K��4D?]m<]n���֡`�-&R�U� �M��IEk���^!h�WQ�	��mY':�m�f�]KX�y��M(����\���n�"���W�B���J�\����c�v�ek��m�޺��0�|�Df%}Y��*�&g\��k��fAG\L(�(���|�p�cQ:q�s�S��@`��a%`9Y]�m���%����S}6r��~dz^�u�o
�\F	��=��ĺ}m�㫩�N&���0����w�?�2�������� �*�8n�������:K�����e���aͽ�R���P���u����~�u��l�P�CG��"����$�c`h�bMg��&��F$\g�Gv����<d��"��y���|�Mb����ͅ��1��Ʋߠ�:5����0�2�۵5���+�Xq�T2������7`��߸M��c��	�j���b����S��׹v>jl0*RP����������l9�Kg@g=�g�aOT2@tH����".
���i4���P�Y�(��`����y"q��tj��/c��t�_:)f����w������4g���u��%hs+��c���'���ZgN�������7�O��[��Ǡ]�3��H�V�0�_�\,aL|p�5�>�n���
	BD9g��v�M}�w�\��wR�N�B��8H��E�]|�3�?�&�ɉ�P�lq���&��p�B(E�cn��Tff��+�䠟�E!\[m��<����-������-�>w��GptC��ۥ%I�ܾ�@��_�YX�NEg�يh��v����Z�6��o�f�x�[�����0���-GIda aI�M4v�2�	��C��Y�^�#��}WEgM�?.l�
�r3p��`F_�g�<�*o�7o����l�s�?� Ϩ�b[q����U�������E4�y��/@���u�T8[I�/貧�B�1�4Fr��bb��r�����x5d*	�B����H��cêH���l�k�2�%J�A��52ׇ_n��w�U�n���y���V�v��7�
�|�jųP6�`��`�Z�U<�4UA��	7��!���EW����l�)!o�]?"TCk�/�>G���A~�2�����T���� ʢ&�UC,@L-�:98Ɔ�^�QrmN�A�z�~m֩���xm��\4����_�;m�l��D7�e�xJ�|��
$L�Z�17±U��z5���;�e����W��}��\(�mr?��+�ebѬ��#���}���4s��=���AVvj[�-2  �.2B#�$��Z�U�H�ߪ1ሧ���-��x8�e|�p�;�W�����6㢍�b��eߢ��s5"�^����j���9o�a���6����|�*�n�G�<���������E���Ȅ'��Jp���2�M�;�H@B����C�Q /�x�7k:�$��.\ �����@���OIu������Q�B�v+����F�d���6o��	���>!�KR;i:֢�W�'z$ "Zz��3�<�k�p���L���L��q��6s����M�9�=D�U�ç�˗��՝��b_�{���Y��Nя�9Z�.���4s�:�)�BZ��ƈ�
^��E��[�Kg�8P4 ��n|�k1*9�����6=51=��K�t��^'Nn?��r��ѝYL6b�Y��߀ґIةR���~��0'"B�R�r�����A���']u=��U�2��)��?�y�E<�����$����"�	,��`̓��D/)��$�%,�ն��d'�pn1��︀��=S?�cMs����g��DJ���JYP�H���7�>w_���!�s��q� �JUY&wVМX��vâ���;�m���E�(vZ}綅�hf��0{a|���3qΩͼ&�Ι��l��e�U+��i��6N�?7��Xk�`- �������m������}���A8;DHu��� ���=�nC��M�	�PZp(�d�ՂN� ��i�U��޻�C?�	XzD��<&��c�c~��*���R{�[����SVݠx��AX��<�P�4
����$k�
͛��jw��'DaΚTa&H��(�<}�P��
!ݥ��{��`שX��Į�^�6;f�F"��5�4��ZR��*��:=��X%RbBWzhP�v�H��d��#"�ض˻���&�����_�OncO	)��ܤ��Q
WǫM���lC��:#O2H٢����Q�Uς��n����q6�m?G���U�n7�g��bla'�z�
��(�Ã^-��vI3B��!c�����Q5��1;M��? �ሄ����g1҃_{��H��Yq�lke=9�������@~}�m&��W���l��g�����S:�_���SOٝ����[V��2�����&���9������7@���"�L��Ҋ+i�EA=�w�OM��Ia�߻��?�,au�Ԛ̡~7D�|�e,�nx?&0�?�pk(��JUd�u����_uRN=������h@���uEU��*wgV1��-�\�z�|<_��/
�:@����'�����k��������x)�Q�;�s�1��C�q��+���-�����gL�N�Y������ѧ��v���}�>w�G:�i~M������\_5n�e��W�m龜ܧ>%�X���M�z����i���8k ��������}�|<ɲWf�-����U��� �o#ڛ��3>�� I���cWp����hs�N�uZB�!����b�) �+��\��T��u��/��@Dƃގz'�TȿC+��w��~�^Vp��76p��9hd1l�<���<�kiNY�:Ԅs�F&�6�됫��- ���ʜ?:2�N�0�x�t��M�)P�H��ݲ�ֲn���D?�X�=���߹�� �}���C��_}ϐ��6vu��Gj�]�[�����}q��s�AL#�k���M0�̀r��Թ�olG��{h\�±�6W��I�����y�Fc�Z�s}��I�:̧���镘�`�F��o3B�9�J1�,\?��sr=!���	�B<�#�Sp��<���0��Ғ4��٠�Y�0Ex4�\<���s�~�]�:��V&�G}����p���Ś�g��w���^���ٯ�z4d^DwK?�R��'��������'�~�TC<O�J�`$#l�W��� 0NɅVn����HE�i�̣��h>O^eÂ��}�1��TI*��s�����=^��ϻ�N���� ���tڇ�r�5U`��U�`4E	�;�� ��	xܜY����ls��,{2��u6���@=��ti�E�(�-I�����I���q#�#�ɻ�q�F�c[S?��[�W�)^��+�i���0H�u�����%����[n�ɽs�y���	��g�|�t�0�d�x��r��*@��������1��_�~�.¬2�]�N&ks�W+�}Ǆ���X��w�3_$��M	�d;B�az�}����4	^�̆r��k��$���;���f�Q���ϧ�.���b�̤469��/Y�qr7�g�_Dm"�<Y���˪��b�e!k��>t�%��*�賗!�A�p|Ԁ'�-��@V�B�h�ࡷ �/TyOol����L��IWR�D �ʛ��b�S��ո�]�]St|�;@@Ix��F3�<���o<�P�[.�K,�{���,��3��v��	�<�x?��|�ٚ���
`���w����3�%]9�R'��b޾r��t��?2�^`���F�_�5���?bC6/F\5⺛��G��n��	�d�W��g�x�"I�}�����	��#�a^���X����ՅQ8���֎����"�>ja�?D�QaW/�y�V�l/z�����XR�H���k&��ЁŃ�r.7�3���=�-+�ߠ��ڦ��ga��]�H�v:>>�0�����*_oOzĔ؁ 'C#4VD&�� ��<K�n>�KJ��S0I��U�ap9�?6�W����φ�!7!�[Ɗ�G����Il�5..��U�Đ�0H�U^��^��lZ(���*?9P1��"ß@$T�z,zE7����c-���yZ3w�[���)���b��H�g����V֜8��l?�� �n�J���Tt���_�������~Y7"�Ҭ<�T-'";�<���[B"���~ߊ@�M!�I% �ъ_.��kWr�Av�y���}�B� �Ov�ڱ@�XI!PO�d���b��^#��h�3���&��Z�V�b�O{�}#�c}K�ix�e�XU�93��󫄰T��qVǺ�����jn�X���^�C�����vY�Pz��GlS#ԾM+tV��5`m��W���<R���D0�9�=�1��P�Ӳ)M���G���;���A����6W��I��&fpH4�,�@7�Z����*�r'� �n`���tDVgu�Eq�����=���B��-)#�2O��m���Oz|���B�ֻ7KeCj�uƅ��8�������/����i��S	��}�_�f��v^n��u+���ا��j�:s��L¡�mӅF ��Ԍ��B��@�G�3���m��6,y�g���L�J|SM�
���F@C�/���V/kob%RX��5>p�[neq/	���I��c��FB$�e:襜g^��Czxn��ɋ�yr�cs�%����q.T�y���>����ͩ�J�M�4�)��+�Dh��Znn��jBvz[��n1�h�D$���R�n����X��R��<�1�+��P �Z
���y���/�9h;�h�v����,$I��}~��'��`3���3�������ɪ�L.�����c~ۓG'��/yPk�� �	�פS7xy�h�&���Ͽ#,���07�%�G��(*�h��exDAuzL�G����+iz[W� �S>؉��[\�Oم8K��������B�T��8�9u��:��"*uXz��i��.R���,"�"��گbH:�ʸ��c��&)Or[b���X�Td��<l���i(���էQ�a�;���(���g^��X%Ɲ�iVL�P������ #BFF��iF�x���W�4r�������|��s|�[��}E'��lX	������/hQ8���?�W���b����m��B�<��#9S��R%:D	����Cw��-�Td�C6݀��)�&V;�`+5`N�b@�C׉̆R��J���\TX_�u�̿�KpUe*�m�&P��>�&9��GR�&;�6_Z�0�a#����tM��x?`	�%A�iL�D�	��,5���H�0)jOJ��S��9K�|�u���S��H�9�U^7�RYF/���7g���$�y�s�u_�>��ƬHh��D<
��ΡX��Km��T�5ʊ�%s -�����|��p��d�.�H� �e��A6'.��@֎����-}�F@�T2R�.�|�I�����{B���R����fR��T��j�w_^Z���O�asM��"F����A��R[K��+���ZA�}����a�f�2�8�z�ɉ7��`/�6*��2h���kTfb�F����Ix٥2��P�b?_cw��%���o����Bq�5|�3�/��#��A�v�EMGA"Q����b�:д$!�KW쭭g���'��`,!I�\�a^�\��k�<�4�9�i!-��s��H�ٓ�]#�҇,���ʆ�'W}�� �D�s���\��u�Z6�a��A�`C�ʌ8�}�_}�=o��a�v����6_���
_/��C�7��u*������Ȁ�?��UN��|ie7�~"��۬�rq
�^& �:C�m���i��f�	fʙ�V֍�z��f�P��U��h���7S�ݼ#����g�7����t�Jew .\F*���������r��,љ�S��.��ƵENѥ�D^�H[�P�>�N�R����7�v�cEc�l���y�jH��<�<t�.�ѭ� �yHHln�����H9��O�=w�Y���Z��b�L&���Ud��qʨhaS��m���03/�� ���s�wHVq�[�dV�:�um*t���&�.A�}c|S����nZ���d\?��'�r�����he��X��$�6E�n���vYʍt��I{E���I$��r���i�H�t*�a%$hI `8r����K8�����KT ��O�<{;�8�mZ�+oU���]������<�߲f������X-��Y�K��Q�^�ξ3�F3 !�&>��H��Z�^h=ץ`���Z;��(���!�`�J�@��rh��\@'_.�=w��_[F)�S.$�y�
-Ɇ���N��0޸��f#""�������T��#�,Hզ�L6U.Ԍ�(�L��l��'q����g�͛�տZ�a�v�nivʑޏ�Ư��q��ņCD���+�B*��v���_8�
p_列%`�E���3LO�8t`4��ŭ4�tsʷjΗ��?�"������V��f�=�5�}ؼfg�un2q��t�j/��7��J��&�{�
I�{}
�r��dtM��m��3Ev�D��՞R��bn��޸��2xJۋ��םS�S� ��#/Wps�&���Hx������s��R/���R� ����R=�nQ<�&ыE�vw�����X��ղ���cnO�8��*)G���J��Z����N%�4��dJ�ZR�ӈi�V��d��MD����h��,y�"��k|D�8�m/ߍ8��-���FԒ����06�ASa�6��p��˥6>7�#6NOd\dq�-�����њ��
*��
L��#�����	�YH�DI���BQ�H�� �i�=��������L�U�cC�	����5���FÉz9zm��t�p?��l�=��j<�Zsn�l3��mt���ဍ��Z����,��<��%�^��'[t�ͫN{�۔�E��K�����]H8���촕t�㪱�{/T%��Z�ΣX�SK�������'ᐟX��M�6^0pi�Rr�HA򤽫����t�ꃫ���0�{�S���B�>}h-�(F����C3A��>�\�n�A�V,JN����?rn����BBv������9z�eo9z��Y3/ƆM� �f�p��{��Y�l����ҋ�\.�b�k`�5Ԡ������q_K�*
!�JP�L����+ʺŒ`�M�Q]�pf �wxmBv+q�t�W�:8�I��ڢCȷ�����%��;�ߣ�^�ȭξw3�0m�T�%Bx�"�o0ϕN�Vv\��Uݞ���']�bV���մJ���>h�l����/�}�{S����?�T;t�p���L�g��c�g?/-�
��!��d ���R+�f���Q���C���C.�ǯۍ������h�rnQ����# Y�#b���P���B&�!Yz �U �
�-��Xab�.
�s���r
��O=)I�����g�!�9F�}� ���1ɀ�,Mc�Ǯ�ޥ�fJ�{�o|����}Jx-�zN����o�1�!3t��p��1gdѕF�tn�8T���ݟ��7؊���^� R��U�;5�B�o�MY�f��/� �<�˲ᓯO�&��\!�ܹ���5�+�ѣ$D���^�_	�t'x;	��z��Q򀙋�:1�ԁ��������r��)�5U�'.�S0�"�k�����S>�}i�ŖZF������Ý��K�I�]����<>x�C�ۃT����u<%[i*+6 ���$��s {�ͣ��W��GDp=$t��_>l�sg�Y�svD	
�*+�\���I�"?|�u�g��+}Ï �|�l���?��	��옐��롚�.���PWYm�쐶n&��Z�u|Y�����J��\e
t�3;K��D�,j�n%{l�)�sa��'i��Oy2x΁����#����ڪI�!^S��Bfi�gw�s�;C��*9��}��ޞ$)JBD�"y{�G��㪰氤���3�5�@J��'�&v�O����!4Qj�7X ]'�6*�^w�7��c���u�W\�U�!�9�Q/���hf�A8u�,u<N
�@}�{(⦜�9eண�(���p�o�k�Y��^���U�聒{3�m-�sCi����x��c_;	�C),;�/�%�g�E����h�(�]���4��f�+��z~���	F�e�Y��������ߏ�\Y�����ƶ�%�m%7�ùa����R���hv�e&ɥ6�R������U��a\���5�m��ri�Q�������x�.��3��[n��7/9�Xd�ܠWޮ�ʋx,�22�����s�4M�~�D��B*��!{y���}C���.�c1�&���M'��5��P n�i���1��R�-,݉tg������#7�O�mxT�������-�D~���C�)Ct�H����LdGy$g}R�\}�yD�Y�N��D�G$�zV�2Ӫ�t�}H`f���1*g��l<�u4�ӂ��O�`9!Բz�8al�&�����&dHb��H_8�5�q�a�ٵ򉏀޾,M� #'9��צE���1��v>�z�Tf~�Y=�DNH'<8�qd�ѱ�]��+��--J�2����Xپ�8	�{&�[E���L��<2��-���5G��� @Ax�>������K���<.���^�%lF��eq��p��?�G���=X2p׿���-C9�zsa����L*蓻O��-F�{�հ?�jJ�����l���%-T�C*�rlE�r�>���7��נJ*�gC.9��V2��APש�hdv����=:���OU��� :��2}��p����;��x��z#���g�9~#�rCL;BB�D0�(RC#yG@1�.��Ծ��k	ō�̬Zc���o4�uG�5�6EU�~[��bL6��]T���k�n�n]GK�rƋ��6u���/�n�Z�p���F�srܕ�Kz�+)��'C@�s!~�k�G]3�nv?I.�p��6s���t�#e"��0V�m~;qr�/jt�ԡ�?G�d�^�Rkf��w��&|Xa�M��~oV��%�r�������-�9G,�n���<�cv��82j�^��ex�Τy�Sf>Ш+q���n�Ȉ��/uD5��~�����Z�˯`d���:�Ox"��cC2&B)>"�&����-����p�(=���#'tpk�@G�h{ :��R���v,?�qQs)�V���L���9���@��7���+6�!;чt$�"h4j�d�K?��:� � Ǚ���lwA������<����:�\ӌs��������`G�"g�Q\�aARJ̹�P��Z�Υ�^h��CWm�	ekU���<� -G�|�K =�L̫KoZ��JJ�|���t�i1d��$Ԧ��o��8R�.��/˦��f$N�!*%P�>���7\1�7�W�W���O�H�"$�b^���l8����Tȧ�xZ�,�2�t��`�ˇ�`�
��]�)��./���Ԅ'���L��'���Z78A���/<���r❫BMI9!���e����� �"q�z�(7O��-�"��d�SI(d���5����v�$=}4�b��.j�*����q:~��J��O�/(�qV�{������ᢻ��:��׸f�US���E��*S �N��~F?�m*B'P��
���] ##9pdwM
����ڰ*yP�C=����B��W��HT.��84���~9"���.ڤ�� 7� D�X�y4�d��"!iR�:70@[���*J�7@�𑢼FD4!*VNfj��d�?���$s�'����� �--�"Y� ��P��\Ho��ɩ��Ga||qG!��E��$F��	j9Ie�E�9_���
�%$� Z��Q�]`��?�A����:���N]<	zQ��^\�dnn��"Ӧ�N�2�u*���yG��t��ܫ���@�4o5O����8��?�s�z�5҉��f�6{;�M����B"�Ә��r�uICxQ������ܾ?:ǫ��g�d�y����x�E0=��e9��~��H���BNp���.�TMk�p:�qQ)pM�;XM�B9(�pZ��%�WG6���}[a��8��������6�E��ciA� V�������m��'8�90�e|�k����?����v��uպ�����e�~pӯ�1����~b*�i������c6�6H��(#3 ���/ߤi���o��	?���u#"4��s������8]���`���ڦa�yv���{�旎RD���7@�{�"��
�.��6���_�1��:	>o>{���a"l���2��0Υ�ڄ��l��26��^=����k{	�[r����m��?)ED���@��# a��'����<��f���e��7!W����<���\���"Ҙ�ȹ��F!&.^!F�~RL&*��I��%�z-Q��E�^�&�I�  ���#��ϸ�Ų=��,���V"T���f���]���šLFI��QRE�҃�T�+z�u�����v]%,�;�Rh�����?_ٴ#��L��~����@�Ku�C��~D)�Z��q`ENG[�����$�k������;�<����?�hw��XL�ޜf�w�j:�_* O�F�� �IZ�j�K�;ٚ�F�R���0z�V�=J\�ą\�*�W���50�/������MN��׿����z��G��T��;{�Ak5��T�*O���#��1V�L�V�ĕ+���j��1b��Q�-�n�1l�!��ѽ,sb.����c3 `����5���fPc,Aer;I$�9�3|��Q�4Kwv������
�:5�h�ӗMַ��xUd�P>3d��v>��wI:�U��֊���T=�)�p�-_2JX��XrhP�q�Ф�Z�hw0xA���'��<e�Ҥ�
~�(�ٌ����k+�$���v	��¤x��mV/����Wd��g�^�W��*:���Tq��f�ڲho���5=
A���Ү�4�(z��8����~Aժ����?��R������P��[�t��ł�WK��ߌ�:����l(1C8yyDF�!%Y	J�Y`�~����OZґ�R�~z�#}��L}Z��\k�H���}*�kR�3�nöltI]5��	��S����x��y��2�uV�~�{z��7�T&<Hǒ8j�Z��%%hAm�%b[��z$[��=+;�5��Le��m������I�L���殙���h����;��7��V�6r�l���j�w����c�{��D���AL���e�Dq-�h�E֭+A{���vў�~$"Nt�B�r�Ƨm�5�o�ܤS��E�QT[�\�Tڡ���4tR	�,�Y���D)�J��J�c������0E&�i$h��@��,��I��u}���U���d���C4�h�M����Y ;�|b~�$�㎬��̋bI��4�����u�m��YQ�{�c��{�e0��F��aF�u@_���u]W�ZM�'[�]Bi�	��\Χ:.� t;�v�Q��ۿ����.T���'���D�Ē��d��2
c�g�i��\�?��$�y�V�G�&-���IX�	�I�R `;��T_9�0`���!ct���E�*LJ�&�����h0V����W�M)E Ng圩D����0S����G,��A|��U�����	����U�(5M�o�̟7Z��[��X���D_��@G �v�p�-7�T�fv�D�������mҦ"VE���ܔ[��b�1�:�t.�鴃���\����j蚄Dh�{��{��ɮ�7�5p�t�f��\Yƣ�F�oR��{�~#(�r��e��4�s�Ȝ�>��,�&~j��>�nc^ˌ	S)��5�ʡ�eI��F��,���S��i�{(yG2��8��Z&�N5e;ޜ7r�#�6M�t�����AiR.Ƞ��+ו|�7�������6�`�"V������9���xބo��,��^C,�뀶�
���J��
���E�4�jmw(�Û��� #�z�4����y�/+��Z��hK8�2�?2Y����f�
�<8�~������7����|�;�#��O����$���Z�M���h���]�p��͝Z)��`0��� ��xD� ~nX#X�XI�U��Q3�ol��,M�`-�^� W*R��� ����|7��lm�Hߖ�7+ٚ!X�(��J2
 ����s������b��Rw�r�0r(2/���p'j���?��\#��R���a*���{�����T�{��d��9K^��-��i����"��Nɠ� �JŢ�eAv�t<@Np��"�z��pI��@/7Pi�,�"�Gޚn��l�N����e��C�=�|g��fs+}���o)蟅e$�)����	�5�w�x��I�B
�+A�W��٬㫺�d��
� �p��k	�t�N4��?�Ɵ}v �eD�������!\�lc�ؤ4�<�#D"O�ӿ@�D$� 6����5�~~7 )�̈́x��
�R��B������V���@�18pC K.!�Ɇ]k�0Bݟ��y�.���+w��Į���'	I/�y��*�����tJ\@G.�ڽX�3��>0�~��,ê0%;�`�swu�ԏ�k��#M�?^��(Q�Ш�>���Yr�ڊ;E��Ǽi�I�%1�>��|���,�&P^���ŀ��aG*]����I�X#��slZ��x;�'P�mo0ƾg�'�Z������U朸u�iS'K^b{��(�B5��}܈R� ��%]����?���M��_�4�j�'�V!�o_��:���:�]������^o���5vY�c���f����5I;�䇇��o���[���b��H0B���B�B�Y֦�/</�F�`p��8��:�i�KƦ$<��F��zڑ���`U�R�dS:��/2.I��BbYSN|e;��K�Ћ,��>�����nMK�e��<b��w��	V�q��cW�MQ?�R��[�m���cy��l}:�!̯5�j�Q�� ����G�*^�&�b�X�"�Dg�J�IBK�oo1	p3�FR�|�R�����#�UV�f*m��=OJ,`XP<�������t0>�����}ջ�S�rCF��4t��#4l�9ldT�V͂�8�\|� ��`����D��������{.4��P�#4l��h��B���=pQ�E�72~�U��*�rH�z����
M�Qa+�\�I]�W�s���+��?�q�|���C����DH��ƀ���?x1�G3X�W8Y�`��̨ W����N��9ϴC��/���"|�P�ӈ�ξ"b���6�b��d��:�ɝ�ك�>�`�D�n<��]'Ax�hٗ�|g.��1�����/�DCWi���a�s"�/��P�;H��v�����蹑o���;���m��Q��9��`����O�5^-M�NJ�P�����sT����_��Ύ����+�)n��ZT8�N����1����wۤ�y�h���`����vC|�@YOEɔ#o[~�hR��7
�D5Դ����� Q��i�����3���H��0�A୫h�1�9��p+� �]��⛦Xj�IR:bH�@M��,�$�O��:�0�$ɘ�a�����#S���N��M�cX���k��n^��o�:�҃��5�FSs��~Nq����U*S%�Bn0
��D0��X��T�l��aDd#�����̧���� �
���+`K��G��]�;%:��SN�c�E>���.����Ĭ�[�^�.ж�֝�q)2u:\��S�F��Z�J�jI�����rdBғw��d�ƣ��w��8�Vc�3��ge��\��x�?L�'`�"�����|�ACƻq���e���s�7�qD]�^jz��=�s:��ɻW���[��i	�5̷C��ɝ���h�*�".BAYIH��j]x�^���U�;��@$d��B�H��%"RG�<9����XIeι1�r����<+<qMN��kA�@>BܣTT� ��f<�F����� a+b-H !�T��>O��d6�+AdD/��ƍϽ�[DRE����>��KL�zQŮy�($�K�N��7<	�'�6��<'d�Z޽��b�уk��-�s^.�ԋ��ǿ:� ϭk�2���m�z=7m���X�^���,U4��Zӿ8�،6I��}	�>-�#�O�$I�Q@�	���+��� ���4����s��������ȳ��j������_<����;^�\���״.������N.���x� !���C��F����	�Tc�O�U�><�8A�������,��H-����Y���P�W��-��j�tW�u����?�E(�6���ұ�@$����ʄ��>:�Y�F𑩓�lU�d�>.��Z�`=�P���+R-�p��V�(��+�O��*�y+^�45��
>1._L��&8��G�[�wi< 3�!$�F���B�:�En��a��xFI�Hv2ӓ��x�:�����<O#�_�82��E�
�"�����'�c��۔��7�X8�:�+��(��dGjO��z��.�!8�������_.����DȀ�Y�M�lt x=*��_�������䟒\$Y�3��,�7�8s��Wl�z>y\��L��
�0u9D����F���,�ŏ��ӛX���kv��'�@�{+�f>b>���p%n�(��E)�2�"S�U.n�5$���Y��R���D��`V+�VB��Z� N��b/�dĉL�l{(���Y�kB��`�\�l��ł�@�a��DӘ���F`�lT��9�����p�[1��d��,���,9�g��6E�ϱ�������b�w�Z���2��͛'NO���ciC0bx+��b����<�Izf���	��|'��9����	�:�ˇ	/=�gM�9i==�;f�mR��2����1���d�R�z�:gt��T*C�}�6�M�t��Z�+���唓�_�$82Vaӥ@@??R aU�m��'*���'a�i��Z\+Uɏ����
�MTxfR�젓�n���;)�/X+���e��^�6��B@��b:���I���}M�Ϙ�i��1�ןs�q�E�t[?$��^���z#�_�g���Z� �q��$)��$(XUIp*t8��Ov�aD�q��甈����9-�m����D��^M�_�NNŬH j���,p��E4Z7�X��`��&����0�RN��}J�p�X�z@H�ځ�����	�Ym�D�)v�+��6�G�<�>��s��Ԥ!*O�>rfܒ�I�^�:|39��jS�R���Sgb�Y��x�FA���	f���2gUe�PP�M�����é! u�dHd/��p0&��G��cT��K�j���D l8��2y蹏�����I\Ì�1B�~Ը���N{�]Q:�Ԥ�UE� *�?�r�^bEL��ZRJ\?�+�&�k��aB�J�?�sD��##1��Z��Hh��Ľ������S����N�%_�W�����RC8�{"��PꢚN9�E��o�o�7��F:�H �Q���<a����@'C\��^~n�H2I��{|�y�[_ou�	��s�8Y�F�{����r�i�Q�1� � �P�HEC���T�����)
#�S�I�I��d�y����2d�2Ƃ)�f-%.�kC@�!����<5D����҆���:����n#�]2�8ӟ��y7�����ަ������f�df��2��S4?[d��-��a�9���*YZ�M4��@��8û��d��j�g�_:^�� ����\����s��J5�%�ij��Kɒ6��{�4�����t"�M��x��;>�X�d��!�}:?��@p�	�KC&}r�섳��t)d,�*M��B���c��?Wx�*�! .�DA�B�y2��F?���]vF�cG$���YAؕ����Fx ����{I�ʍ����������A�i~UA�|Y+��j,-򏈈8�x|�$�ʲL����D�p�-�2���rē����FB#K�y^4�N��MqM興�	���E$�*�ђ���a�r8��P��F�&���in<�h���ߔEi@=4�6�Gc~ߌ���n�e~���R�\�0��X�KHaSjD�Z֠s��ӲF����^7eF���>���^��~�y<����a�w��tU��� �Ia
",�W,�wpRB�@"�CR[�#?RKiv�O����?nr��6�C�'�z��y[;����P���h����{H��M��Ϳ�t�$H�c�_���J�{H��ϟ��;�������w�Lj��R����58.�7A�>^�I���ӷ�{�׮;/��e�G���qj�͸���R��"A:>�PY�cZP���s0��ZW��4����O���#9��X��ڤ���-�˾�4�u���8}@4�i�КP��>g�g�7�ț�4\/»�9����@�('c�����I~���8&L�.y�;JJ m�sģK>85'H1i�=�u95#7I���J���dE
U؈��,y����{E�ZE|tT����]�jS��|�*Tv�^4�4)A����j$G������uڕ�nێ���'�lK��^i	OU�Mu#@�헶ē��P��'I<+S4^qo\_ 3L��=�.��l��o��D�n�=SЫ������ݗ!�G��Y~!h{A��w�h��}<�����$�"Tx|���;~�E,�t��J;$��^�N�M�$�;"�I�ZɈ�s�c�`�s~�b��g�Y����f�����tz�k��������,�8�D6i-�k�#%�+�
�@�,��cA��\T��q��5�#�9]L 8BD|;i<z6u���
D���F"E�}��;��B��^�Nf#CL���#T�^�N�	�!w�h�Mov��K��i�CM��T3D�ݒ���@X"đ+�m��2�D�-�暖��(c�����η�Kw�_�	���,A�YI`�}�S߉��Φ�������I����xA����]'t�|���{��������o��V��q��ήr\���������8�8v�9�'ܭG�����5������9�m'�����n-6��r�`<Ρ����A����uM��vY�S}�3�+n���7^��m1��p;m���Y`0EƔ�c�|O�\�@�&��1��Rq������ƾ_C������p["�?��ӵ$�<݈�rM�1ʍ��c�lᚻB�0��#<����f���EK����lӒ�9�m���t���>�� �����,"#iG����5��l�LY���?�cCt�C	��g���U]�RȨp{� =��������p�J�����.���CAy߫�ڑIsn�A�s-��׺M��e���F@l�H�x��z���Ӏ�Ǎ/�M5�,alƝr���7�K	ް5=����8�a/��֔����w����n� ����y��܍����#"�4fn�듎0�(�5'��v]�)��M�F����pA�f�G�l�Y^��y�4���*�"�>d����LV���m�5���2ڴ����C1���]Ag��|ڕyFA�A���U��p��=�a��3���\�Bp�U�٧N���`�w�5`��ƶ8����� \D��.j../�Ii��I7��|�y}�R�z���k���s�Ӟ��_�yA^�;`��'�%�sT珥B0�%�a~�3�u7�6��L��#4�o$�$�.]ߵ1~��Dɝ`R.�%(����rG�B�q��̵�"fM�s0\?#~�K����l��5;n^��S!�����]�g��=��q:@Qlwr��ʟ����1����!���f!�_���(��ݹ�<b�H�1��I�ׄ���G��΃��X1"�9�ry�͵�TyR~n
�S��T�*���5��R�?.���M~��IZ��b��)2��M�Jq�O�O���R*���Bw��yߗ>7��@��:C���b��t?����sy��R�9�L��sɹ^$�}�B�iS)E�<c��a��Ra�W͕>_��}�[�^��z�Sni�꒏�WU�uۨH9c%�Oi�]�OnӷĤ �+���d��D�j�f�5E�4��(x݆l�ѫ��I���N�8 �'��"N7:��BG����D?t;g��hR�mD� �Gs=Ł��8K舌B-���_cɲ�X��t2lj��kpB��!�P�4u�l�n��غ c̦��PA�M�"�,�5'�@���Ǭ�*n&�˅�	� �	��!�[rV��xы�`�)�[�0��� A��m��ј-�Ƃ-L�FC�Dg��M�Z��u�U����.���z�B����M}�<(�����7�5w��x�(KBB���ǧjS�����Z��K\,�^D�&
O��v/��U������\I�a���E͞ֈ����0>6�% �Z^ .�]c9�gM����� E��vpp.9Z,�R�u�M��I�=Ή6}E��p�ɇ��p4E�[�6���t-��ϻ�Y�F9B)�z�	|��O�_�)1Kf
��Xq~�\�D=:-;��* 2<W��H
���a�z���Z�dI��ln�K���c����y�I۫ΟX��M���m���-��p$�^�M���p׷��.B�j7D��F�:8Ph�G��☾%TPN�A	��2D���poW�b��i��xSz"ύ4~Dĉ����G��NK	i��e���7���^ .זt~W�X�S���y=�:�����*�&��=��4J>��e������o��G`�5����9"i�3�?+�F�1���.Ѻ>�
�WR���g��VT܍���6�*G㈲����(HY�"pY�&�걨��Y�u$D���Eo�z�G7X�L�F`�&�椥(��d,�<�'Nc���[��������)�H�"�R>�>���m�;�r�G���~�� ��/�Ʋ�%-!]�}�~Ԫs����C��B�T3��4�`R��a2��Դv5!�|Pf�vuF��U�od0-�}�fO�?���(�YL�3�å?�����H, `�&�N���1���3�@;�mQ�S��r�����Q@<���[8-�9��J�U6��)����d��f���x�t$#���ܕ�6:Q��{yT��4[�MH������F�B�
#�j�"d�2c�JZ���^F���LN��MjH�0�]ԭz!t[�>�tq^Ofu�b=G����)@0��^�=�Ρ��^�u&��V I���T���27)>Bu�8�8b�$#A����`�E�^���U�şϿ�����:�3i�Q"��5]T���|��%��L��P.���2�*6
�
�S�ND"'x�Ҭ���7 ���p�/!Kz��=$+N�xޱ��8k�V�HL�:"YJqR�zEz����skX9=�_�t+a=���/'�54\���F�!��H4d�aϤ}T%��wJ3�kjG�Zs}GV�t*~.7�ױ7n=�;�c4�4����M�cN*
�́����¸m�o>��1����B�/��0�.5�}<���F�<�	�h��H S�����g�kX(Q��g�������X���5��ϵ|�[�h���>�5�ae�#�8J��:���D`.^ـ�(�S<�>�����b�U�n"�:�zt�^� ��~�ǩ��ǣ]��%��5�!~2)��j�O`�7�~�]SaU�;�Ĺ�"��Z4�ܩ�>�mD.�ut)b7���2T��L:�B���b��"EY"�����%�_��;p���D��݉1n[/0F������JUrA"!	�}��w���$���p�����m����ZH4h����]�t\��H��8R��\`�;��f�v�j�U(�A���>�rq��'����w៿ن����C<=4�kK�
&�SX��?�Q=�g�5�'nͤ]�ߧs���{ӐS�G�`�?�ex�����}w�OL$ ʒC +� @bX��%��帄O>�
��!/^�w�{�{�U3<��ē�>
��￁�}��r��E��E=PD1="�È��l.5����L^m�y/���s��|�������`ͫ�V���jB�׫j>N(7��$�C��{�D:(�B#�P�{|kw�{ڋ��Fb�k�q�X��r�Ex�;�IN��m�K�MT01�$	�5�H�[{mC��^���w߃��3$)=f��E�q,�TO@��R�
H4�����w�|^{�M��rߗ_����F��y�����@��$�~-]b�L+�w/��"��c��ƽ�L]��n�|Hc��9_�H>^������5�7�L����0����_�BIiv:��b����'��Z�������7�ǞRW�8�Cj�~�w�x2xXZ����1����v���)�O�x�����{������!-�x��c�V\�AM��N�����kvU�����������ex�-8�9���CP��_�����oކ_���o(S�k}@f�P�r�c�z�i�<�bg�����!'�UImݠS��4��*�e޺�Z���i�r���p>�}��qBY�|v��}?F@�)T�>7�8��=��~#�dh�{56��>��������>�ׯ�H߀�h�����N�,!K���~y�ᔮ��Vh��(��.���������bs�D+�TrJ����~��K��W��B�����o�hr>���Rp#>�ɥ���(�@#1�����us��}Ya-��C�u�|J}n�l�c��w��{H�/m��Ǒ���W��/���G0�܇Oۤ�"�����A��c����]������v���������n� _~�1L�U��7����������{�܀�G
ɥ6M������3�f�2�/&����$̽�Hݪ̉F|C5�xVՅ�A<v��9�SLDDđ��G���;Rf���� +}	?z�e����E�Rs34�bo@ELߣt�﾿	{��P]�
����3��M���4Bp�������b2W�`#��!ف7_�ÿ������6���u?{/��]����è����� �#qہ�����;�A��>�7n!�t��D��{k��/߅������!�w�.�<�I`�d� gs0�
��tr�ߛ@��[o^���
��݆�`.]���#�~�4�߿�����˰�h�����/?�7��)llm����@�9b��9e#""���}a�g�N�'
2t�% %,R.9����<Ӏ6��BP��؋N��h$�t w�G��g�í[��ʅ�py���so[?R�k�����!���Y0w�z���c�o)�7�x��|�ۛw@�}x����W�"<�ï��H�e���4�NYБΠ�+����"i�r�_��W�6�t9㈈�\�Sx�z����h�ܸ}�נ�� ��^��q������G��a4- ��9ͣ��p��o\�_����!�|	��<F�����|��擥��4�q,��bu|M��z=����?\ؼ�Ι��+�p��B�p�pn�h��}>Vm��R淮R�"�Ij�Tϩ���F�yY�ለS��'e��z��P����⸚���J�a1�O��_Oa�&���5�h�WhDM�� ��Ԝ�N��2��=�4�HA��5gbi�Dr]�f��������������!\L�o��G�㷮r�j����+.����p�"�/~~����BI5��Ye�����M/	bum$������&��C�	�R\*OG�w���^ jy3�֜ڨ�PD�_����y�sȑ:�Ø:�S�Q����M�������>��Mx��E��7ޅ+=��>��^�D���Bz�u����ֽmI5�����ۉ��xb�Z�5��g�ɝ��uUU��+<�i2���w���#��st�ED�����~�8��!ꖭj�ۭ��(yvqA2���@���r�di땯5�{$�Nt�#ſ>��f1�B�ܨ�8L��D�\I�)��8�_�B^�����
��ס�'���'�M�����`kcW64����;�������~�i�ƀ�������5���K���!��+|N�W���Go_����&xN��߱�Tf=����߸�|7��,���{H��\�3���e<' ��8�s�?$��{{��.����dI]@���՗^��:�{����y���ԏ������x<�J�11zpC�:&�FDD�B��D������@]�Q�dpy�B��F���[o���o��
������D��!.Sij�&a��ZI�W"1���ȶ����u0l�ں"r�4�БSHk4�����/�_��M��+�ݾ���aO̍�? �8���ڄ}��`����밃�G7v���!��\_�{�P���HO��!gT�O�B���T�]�(�ᅫ �o��/���8�YIj��5�Fp��^�z�����o?����f�����p��>��~n�ޅ�
)cM�5��?~
/�߁��\��W. �T�7)a����o���-ҫ�O�K��|DDD��q�F�~��8�z��6��QL�D1�6���7ڟ�&��@���!�tH�s:E����/���/@2:���n�<���)JZU+�ԝ�S�y;e_�=l�*��6�+Eb��{�*�8�+��U�{}���ª32|cr��d6�~����w.� ��'`pi�N���@&/���Ar$��������0�|����.�ε>�ʤ�RO
�u'g��W`�^����ݘ���N�ﲜB�$-#���P!|��7�7� ����`kc�Uy��Pz��\�E��O�n|�7� �ޠ�	�x�:��o��x� ߺ�%袆�d�}}~��U���@Y$�\������ۯ��e�gC�"9�(B�(*s�m�����Q��}fȽTfNT��ٳ��'y=NLBF��X���v��(��r��Z��[��<�9n͆��p5*��lߒ�K�R��R>,i9+]C���=sD]��bW�s{�zu,��x��=~T�q�̎S�&\߰$��<���&����F�mo�G_|�w�q��Ԕ6{n�H�� y��RB�V���	���w��}�2����ũXV��^w�{��y�R�=B�
��6�������K�����C<�eol􁴔7��=���0�;@2�	��u���psg�	�W�3=����6�Cd4�ښ8jZH�'���x��b����>�|+�#s�gF����ΰ���U��/���%�Y� ��|�����㦝����$�(�״��4D2Ai�������M���C���!l!1�6�h�����`�D���6�H.�=� ��1n�R<����{��/�4�q_�|^�TH$�����&��2��"�!��n�ֲkS��"�&d�*���6�`A���ث�0"��6�睿�Y
W$�׆��¥m-���ÿ�7�k7l�1!�)��=��M4*Jf�g$bQ��O�j��ՃWoB~�%$%c����e��#�X���:���34���F��S��������=���}�k�ٙ� rc�\@�6F��x�5���^{�5��_�^}�((�Q&/p��fB!�gby��E�S�)sh�B�������G���G7aJ�	�Pn�L�؞���H���a��q�Y�qH&!�|(#}L=6�}��6�W_�M����c�?���y�D��4	��+���߄݃�9�q��	�C���,󣶍!S$%pg����1���hL�`J�X�sJ�C�Ǒ�eQ�3z�"����R?i0Q^g�%12�8v�.�m���y�S�Y"'-�Dq&A�!y��f�Q���݃1��W���6����Bָ\UU�w[���(��4�VP��T��?v�K���zܨ�_�9@#�8:H�U��ks���Yp~���G�)�N��%0�C��>ܸ[��TB�&���=�S�j	���4�{�m�������ʠ�s��Q���K,��Q�z���؞�QwV4,�OWʖ8��G>��:���� xlE!��n���\�D���z"�cG�W�Q!7LC68.Imn ۣ
���c{���'H&���� )P�>�ګ����M�r%��oN��lá�A	}�u����Sggu��EDD��i쓐e��#�6��湈�g.�u��O/g	n����[�H Tń�TS��2(��RR�C���'c��&�����-�HJȈ��q������[�RCy��|��^%&i	��x�����w�[dS����
��d������,#.����y��ӏU
�j E��Ժ��d�jGV���h�n�����E$��ǲ��#՜zfkn�՜t׬7 Uи)�˯��w7+�euq)�2��MȟJQ%�궅d�y�q����I��6���>=<HjѨP�7��x�q[�|y��u�I��D�A!@�_ b�.��tu6�K-��ѩ�'B@�&���/y�H#=MW����"������� I�0�c�IC$ ��*i/�i5�.�4S+�~E5 i]��h��a<: U��#�����S��t)����������WQ�9Lт��E��K^\%3P=��5����two�4�Ӌ�>L�n��_{��ퟒ���'CH�z���qa���.�S����b��i9�������3�p$~G�.�u�9؂)���=|9�t��̡��~F���Y�6��s�O�y��}��s�Gj���_�ip����^�x\��rtȽ�2����S��N��C+�L�q����.�@19��h
<_c$2�L�z��66��o 	ı�o�v�$d�rO����r}(�����{�K���)�}�V""N/��3-By<����X�|N=qD�c��8�@�%���8�a<�U�[qQmB���CH��`���w��7��������mH��H`��C���hU0*j(+W��/��\y�eH������ˎ�h��G��=��$�G��wf�sݐ�'!θ�J/�nH� ��'��R�P>�wo}���38�y��2er��t5�Ǫ���Y���^������k����o����j�C#�ҷ*(�%,P��m�Ǽ��IR����ɇD��[S/(-�8�4�T����'��c! ϶@�PH�D]���dH�&������0>x ;{�`zp�hj<w�C�&��!՗HH 5���/�W_z��eغ��K�߸��?�ǘ�C9�
��N�W�dM�Z)�`��>�������D,�rC�GpC"ϟr�lG�DD<S8��|5%r|�hD�{ �Lm�����i�?�۷��Ç�@�n�&yUK�x�����U	��\� ������K�����W_�������å�+p����u�Mo��t�I�U q
%��@j�C�x������DO���!W;���ܽy���Tx��|^�un
�E*���5ԠN�wa��L�����!۸
�����y�u&#�ŗ���h��0��[R$��5�3�X)�;e��)p�tj@�.��S�9����?�i�i��tR@.)�� 	}:ށ��7��7����o���oA+<j�Dp0�3��l>��e/��U��)}� F�)�:��߂���l\{	�Ǚ�u�9����]N��H\@%F�g!<�c+""b9��~
��ӌ�냍x68	,��iVL�u��jY�qҗ���L�|��}8��=<�j�r(ࢬ�ʅ�q��)e���1��p5�Äs�'�
�;�ý;7`BZ�h�Bv	.��Sx�O/��L�`*Ճd0.u`�tG�Ʋ"��|�Ъ�y=@�=?�s��B�a��އ{�~�����MH�=��\�:`r�&��R4N+M��k�0��F�X��[�x��x��$��q��/�O���«?�k\~y��SX��pm9\��f+*�Q�yVXk��������4��f]�'j�t	Y=�^�?|�{����>8x�F�jHz9���k�6���$�&]8�s�Xyj��U�z�w�ǯ����x.��&$[/���kPP]~g\�^ِx�䛛� |'"�y���X�{�<���@�d����>��]���y>b���ot����~J%�G:^���V�$��yĔ#-�/=����ii����*B�5$�`��ؽ�1l���}H�x�9l2��!���s��k%JU�0i����\��B�ҭ��L&��Fm��x| {�~�;�|�'��O�^z��,���&*��b]��i� yS�M:�b8f�>��W��S֝w�N�1�"4�����T��d���wP��·����l�Cغ�D.؂i<�Y�����$���XB):=4jk�S�D�@"R�����!�;7��۟�ï?�������� ����	�}$�ʸ�����*+��.E��gh	�C2:�"�F!N�b�Z5l����00ĕ��!�������{�n~�_s���\��p8�k?g���>�m	�j�n��|�ܛT�X��4�5M!/��8N�lހ����~�_}^�o���q
X�c|��JH9�Dy�Yw�HX.G��XD�����ku0f�Xd�Vh\�r��-��=�u# ,�'!]�8��O��hK/9��K�}6j=��6��k4�{��H������ܿ�O����ڐ�9�u�<�� )���{���d��������	\�@/�����34n����ۇ�Ow�s4p'{���~�$����[���e��ς0�yqs���@�YS% u�%l&S����� ݆l� ��m����>/m
�mWG^�乹�e+�L�3#�7H�?���^f0��4�a:��'�����_���ʏ��n� {�Ȭ�������T"��:�ȥ�R�귑I��`Ńo�΍��?��P߿��R$|[�>����|�XS�FE�f���� ߀
�IU�����s:�&ϋ�
a��+�K�tm��)�!��������ۻ���O`x�E&�ʦ�M+``��^��q�H�;�(>�U �/��)�y]B�M���L���"N�������
�?�@�G�܂�;÷���!ٻ��佭ј*Ѹ�P��� �MͺJ*�E�'I�p!��6=A(�Q�Ɣ�ᚥ)�V��us#�<S0�j��4��}��ڇ��}x�W�#���HBRH�9NNJ)r�l{~�:υ(أ.���{P�݄��?a��p5�>�S��K�zhЦi����5�dO�"��!Ͳ�#�%�G�4�IN�Ї0y�5|���v�8~�������X��ϗ5�eC|N?B��r����;�[%H�r<�څj�����7���_p ܇4���Z�&��ͅ��X����;6����yf��4TF*Y��A�HD���8�g9�~G����/�wo��?߆�~�K\���9���&��eӿEs���F�눈�XE@��t�d��L�"����G$ �d�ը�P�p?�@6݁ݛ��_�6�{p񂆞����x�^ʞSIv���HѶ�?�����d��R,��s�⒱K�����
�g�&#����G�����h<o���w��U��������'=N!��l�
�*$��=�<��)|����!��z�|ite�$M�N=C>R$DDʪ�O�y��.�U1#�9
<oI���������������󺉧�����g08��Y�`�@�đ:k�I}��k����~�k|�O	$u�a��~�c+���$������>-8�
eR|sS���٤?��E��h�z=o��@$��S�}x�}�kv:���%l]~�Zຍ�C�NѶg7�� 1�1K	H���4M�>]'��o؏ӧ�d]���#��������KMMGPc"���7Uo��r\?��W�Mw��#��q��8M0y�
zyF�N�J�Gpx�3������m��MЀQ�	S�'� 2��~o�C�P��i!�
��P6a�n�(M`2�p���7��7i#��:�����h�"1O�A5|�����'޸��]�Uփ	�)H9�fF�}��������ݾ��Ģ��Vx|�6���� ';�����/��o
/lj��ϸ7ͅ�H��DH*!ˍaK����9�����DP�WEGj4X�c������h.�}л%����͝�����+\��:�
6l�H�����VC��9�r˹� >�(F}p /m\�ݯ>����?���1yy��1����I�ҭ�9%/jH����x�s��KS�N�+a��s����h�7C���k��ˉ��0Ox/e1F��	�._�W.]�
m�}�%���Vyΐ��ֱ>��x�{]<��Y�Q:u��9m�Xy�8���g	���!"�T��ɋ��!��KH ~�%|���
��6�����)J�lԚ�2nK �(�	���yuɘ��9z��T%Hh��q��A�	:�Hr(�ڐ�q�z�|����C���~��D���j&95�F��G��ۀ=	��:��Ppp������t��|)�QA�BSTL�ǇD5�W�����JQ(�MQ(�� r�I!��"=e5e�CFq�j��`x	��d���!�r������5x���{�e��Az�W��Y�3)��~�u�����p�����g<��o��wa��xe.�W�Z2��C��B�q��sI)�$�c�7�M�J��H��5ե��j<5����X�q��vo����z�!�_�9L�?�tI[�a�GDD�b��cB���X��l/����jDĐm
�{/"�Ԁ�� 4\E�����z�{�?bk@E˚�z2p���M��R_�ī�=캬��c�#) {��l蒬h��*Y�\�6�(ȑ�.��27�����;)�C�P�g����O77�b�
���� C#�<G4���&�~��/~����L���N �WM�:=�<�9[{�"G�"������΀��Bebm["$d�R�+��p}��"[�n��p������7~��M�&��d�/��"!�5���{8Z5^*�ƕP�w��?������'��e��>��l8�Ϲ^�S�j#��-�p�#��StĐ��Xv�z=��2���}UR��	sR��&G���;p󏿅w.^�tS�3$2y�&�ڤ�5 �	�1���|�~=��Mh>�1_�>"���Tƺ+�1��� �"�&(�>��`��W���
. yH�=�J	6|�d��>�z���T���AE�^S�R������sѳ����Q44�8��P�j���2�h,��]S��@q��ҹ��C��!���Cغ�/�E*��b�.DR��Y��%0������j
�� n}�G����Rv W/�`�)��C��ؐ5�n\'��R���N���V�:z�R�|T�)���|�y�T:��k�[���EC9��X0��������˯�`�e(HBX�F�I�Ӆ�:n:u"�䱌�����J�{�>�/`��O��������D!A@�#q���TvnL|�l�A��k�*��As��rF�����k$�4�ro���`0d�3���8�`<����_���?�+?� u�jpXS[���m�2x�Z�9'� ��XΎI��;�
�
��J��g��*:��XJ@�6���������W�P�ӄ�@]������GI���ř�������c%���-#�����$tS3"��S��@��E�ts��鈈'u'��Ӥgv�NL4CS�9��(E�z���f����5�l|֬X%ب�RA-E:�z���H��)S��)���p�$Z��*=�Ř�%�'`�b�AU�d���s���� r4lq�׋�ӣG0��L|7.C6��p���^+��']����AYr��]���ڐ:�I�p����W[�	c$��B����j[Y	�	���YICN
Vd�q2"�#~��E@�|�j�� Y!	�KϨc����+��@IM���@u�[�h������7�'h�{�y�I��J�jUuuuMOϾޝ}����;�f���T�D�g^q�3����f&�L��%#<��i?;�:�^}���������N��˹�l������a��������5]k7i�� !XF�j��i�����������wX=�+�zi����=2��6�yE�@7;�Ţ�>7��H#�A���V����}��^;��:ȿ���/��o#XTC�!���`W���G ����K���������?���c��l
�nu����zN��}Ү�ϕ� ��2>v�=�hm�	�j�0���-)�t���C�:��o�)�x�b���.�����]����pr�d7N~WI�4��Td��R(g��U��d�s��������Sߦ�t"�|2��\DR�s�g?��� ��9��H&�0�� ���}:���h:5�߷̏R5p�69ڲX��&J���5!���
�j��h�eبÅ2B��Y�~?�����{�xgǘu}�����5j'_�O��2L�SblG��05��1���1�9�?��dü;����N��-1��*�hV�pHF�=�>s��D&W��J���l�W?�O�o�w�S3���\F�T��w�w����
�x�yY�������8{i8����t��Tz�?�� 4������O�J��8��TJ�����֋�`�~NsL23�f�p��;ع��R^.���ǖ��q��y��DtA�����F
'�#�b��zYsD���6��.��]�o�&V�BCWs�,{^�0�%�:T$�^��X��Cx��6�Hb�aԜ���TR�8�J^���f��3�> ���ݦ���G|>O �˚�컁�,��62L#È<{��<�wPs�L�����6� �p���L���0�N��!٣g�PJn�b��rY�eIk���Jq�<jrm�a	����� u�#<���_��~u�0�SX��7���~�`/C=Hq?��x�ӟA��0��D<�Y�#��W.����ן��f����D�!�a��ҳ��~ ��lN���ʱ��� Y���'�	���7�?����0��-��2���.8�߄����:*I��&#X<���ӿ��� i3������X����t�Q3�,��/Hh���C�C ����
C��>���4�٠aRg�
h8C\��O����px�F�w����n͐�O���-]J��^k������6Y]��]@y�8��m��=���ak�n$uhb�s���fy䣠 V@���ޠ�|�r ͢�����1��kr:��ʰS֡X�t��~��p��ƴ^�,q�o�[�����|�֬�) BL
�4)yn�c�k90�
�?f��9|���w��/aE���v��fJ(a_���N�?�}��1�B�i*�0 ��Q���q2�&:�@�����F"�`��tj��F���=�a�Q�>��ԧ��
��3�Qv�bi���p��0��~�������������*�O�γ%����H���O�ЧB"�2}3�aV��[�>#K�D���B0((�� D!�ٜ��"͓�W�	�0�F�R��g�o>)g�(E(\�>D@�7Vp<{��+�=z�d�B �f� �r>���-uP�Ϋ\��/�MmS 庛m����}ضΔJ�n�i��;W�d[As��D]ު�i���{3�����u�Ǧ���(�[��%I8>ӌ{�:���8y�-��0+�ZZI���2Og���`A<�2?��&�y���C@�]��dn����C��y% \��C�ό�-΄�B�N@p�ud׮(����� �b�2r6�9\����@��J40�3;}�ajq�EN��I�-@a��� 'f�j�D`R�D�d��I��rF��Z\בA�2�h���Y����0�N`6;�2��	�z�5�z�w�� ��ʙP����ɷ%����9mHsx�䯰x�Լ��b{�=�I����2����5^��j�k�`�Z��1t��X,�ogwה5���-jo/����9,�ZώI��Z.ʳU����"L��/`��)�pt۔4��<n�]l3��)^��7<���^8~�T{}���U	r�w�L/�|U	ڮ"/�ۦu5 
65y� ���wD8s��E�"s"2y�6��7{}���]�� T�	v��2t�d�%J�1��qU.��D@��0��#�@��f�6��8$@��s��M� ;2Hlze�#�u�Nv��lI�]�nԾ
���L�u,�d5�d~
��װ�*Ȅ�����Q��&�g�;{���1e����O��n�儰m� ���,���<x�d�uzG�k�|��(�AS;�£t��ZԬP�,�|��X�H���������y�f'�`� � ��F�rkl0��r_���fʗ��7`�=8����8�1?�:�jA-R���c(j�tNڏ<o�W��pOs�%w� �N����r6����K��@���3�����V�-miK[�����/ �I����C�n.�1���|���ɉ|uNa]�J���5CD���@��4��D�ȕ�Uχc(�5�A�A2�H�Y*�^+u�N��Q�<�̯Jk6BLU�Y�sbh�d���,�����������f���g�1���ӟ���+8�#���&#���7��}"3���/H�/��%�����?i�V��Hi��Xf���
5�d
D�a쯁�%9�G��LYB���٪�i>h�r ��(��y������!��*�ع���Ԡ�s�4�A�P�a��K
��6�2���9�R�O��-��� �"�;$Ԫ�w��2ۜ>>=���Ff-(1���W
���!liK[�R�@��ܯ�� ��6"��:K��l�׹�]>��I]\�kY�.(a0 �z�(C2f2�Kø�Y�svu@&�����|P2;�W��y$(�Uf� ��E��Rr�3��M`����:�
���j�,��4͚JI�/�Y����pR'�<m��nzMf=Xb�Wq~��aP�<G[�Q��a0�bUi2��eM�֜�Nf�_hv��@�p�Lh�32��霘l"���۩�^{}N�h1[��p��aF8&�30��k0��R�p�k��\R���5�wd ��f�䛃Yɥ�E�]�rE�9q'H����j�Ѽ�"8�IGeօ>Tn�q��:X����%�W��q�:}9�ي�^��O[��-]=)�O�r{lJ�w���jS��� $V�^6]6�`)�U���a5Yyؘ�62�j����B��K��b_Vg6m�gtz�I���y��?�M�_���"�X;E>>A����а�M�xC{�מ~�GJw?��ݲh�����I�Wϒ١)�>X¢���W�(ҍ0+ɢ�[3*Ypns�`D���V2���
�<7LeC7�Sn}0�y��dF�aQ�>̆v>�6��aN���%tEa���!DF�������c8;�`���n���$f�}f�sc�'��.�;��3��3�A�(���G91�(��8( �VU���U�URse�p:�@��%�ò��n�A�Ϳ�����{pz��O^����ሲ�K=��y��1��x���(~���9�;n
�U����xf�ӫ'Oh�����,0rj�un_�l~Fe�&X�1�����ʙ���}8v9]V�
L���Z�1D��d<��K&�V�X��!���,��8^��6e���8ڣ��5 B�$����$?0�M�wӨ�7�����lv�:�\�/��'�9�p��I,�a|����|p���]x���Հ\#yӖ�6�k��^��]FAa�x[&V}�&R���pl @4��
N�������h�y��C� ޷��CL�l6#f�4�9��~T+�z^֎̬%�|x�� !�Ą�H��$W�h~OF�a�כ�m�����3mhI�<�j�l?�v�v�-��@#
F�}��ggg�y5��%2DB�u�=Q8�~g��t�ӱ���e�W�&��Pלw
C�sb3�C��B\fB?53�h>���>��/���B(c�S�]��8(�1F�����k˺	��S�n���yxn�3
f�\���т��}�,�Ra�	���R����<)��c��-mJu�S���^���B�7;��[ ����ed~���O�=� ]��*��2��.�� re��ӝ),�`���K�ǅ�%Gf�-*^��v�# s��e�}Ё�ۯ����$eS�ec��B6�X�t�E+�	�K���E_��2�HTVKa��P!e-a�֡#(���r�?���L��pZ&Y�L����5/E^�H/���� 3�O菞C����:3�.0b���jߏ�A��@ E�*�J�����񎀎�����<T���d�f����tf��j�b-�?�X:\�O2�t�*�9���#�s�&6P[�営��J��m����2~�:�����	q�Ln.[E�f&���҅U��i8ˆ��`i��d25�֬�y���3#Cv�.�;�sO$V%s�Ab�<�hfl9�3e,��b˜9�Ld��dE&j�����&2�~�b$��QY�ʀ�\#�ˑI��(bx-1��f@sԱo���I�'����,���'�[�$�L eURJ4�+��E��G��n�uio��xS�����[�?Nh"���|pЬ1���3�#��s���R��_q� )d���{��6�<�;�;_!
Eo��F�O������-miKM� ncѼ!�9�o��q>l~�L��"�*��i�x�̍tv����$&�R�ZA�B\�}��6#��#��\&5�Ö�(�d��Eæ��MǺ���J�Y�G3�'��3:���E%1מ�bE�y��@��^r�|9x~s�V���-�˶	�*�3�����	h�9�Y�Йr 7��h�4�䋃�j��lg ���6�GD��l�c�0g���5noo���g�
L��}�������sÜU��P��		1�/����K����r��JJn7�;4 ���!����M�'���i8�0�68 �C�`5����C�QC$�)�}lw&������A ����P���
�"0���b�ԡ�Vf�L���0�݃l<���p�[�Җ.�|m$�S���>�}L�j@��C��U5����\�YnŪ�-m齣ʷÙX���N�LEdV��a��UhLk4�ǃ�:�^���u��Ru?�3JȐ�T؜��ه�<���8��D��	�|D�u-o�l$&�G	"���ǁ9��8����CD ���?s>�H$}���?�&5�[�ڱ݂[,�d���)�}� �>|��.,9z�{bO]h���|��C��o�I������Z"	�Ѵ�b�@�A�V۔9�2��4(>8���9�����D�^X��I3���1�O�/����7{nmiK[�m}@.�8�s���@��䖶�>qT@H[!���̴3�P6� /UKR}me޵fP}�)?�$����1�˦Y�x�����ωa֖Ȇ0�݇��9�M ����
���aB�;;�@	�a6I��8�J�3a�&U6�.��'T���F�?l{�L�R8dh�ϭ� �����$�'�������3�v_�&{{��/a<ك��7�, y�b��b�=wt�#lt�p̢b�}Rj��0턦j%E�bɧ7�8�]��bUiD����|~:�=�9�'�Ѡ9�����-�0�fW'�e�+��>�߅��Ԁ�!H�ߣ��(�fϯ-miKoN�dB�RY;^�IQm4~���Q%��-��*�,)�q���̧��1�lI�5(̨v����P�v��Ϫ��!�T�$��pnC�教'-DƉ��i3�`2�8�oIٶK����1څ��m��QD�\x��'�#�"�r<�h��t_{�L_�s��
&��ϝY&��A54�0nG��}��?h&7���. �W/E��*��h��S_
�1�m������de��I��7���d�;T�=���I.Y�����u�Gpl��G��\A���!�g<�g�>�������&NZ��Z��ΚD�d�����~R�f��̧�d
K1 5����
��@�zϝ-} hJ��kj�8�y\B[^V�-׼6���5�k�{��.��w��T,���L���K�-)���|j.�m������/�G%���a\��9����Ƹ���<5!S��g�����`����ػ����01�#�Di�Y�3fA���/+ ���߁� ��)۳K�����u�Q�|�@�M:�(͵����'$�}u�Ҝ�YG��0e�C8z��a�va��]��֬뽞��v��ҟ5(9��(��y�+x��`���`6B��0��^�!����Ii����	�"���Z!m3�/�����o �@f���X��t׮��>0�y{����E�x���l�ǟ���������!?�ΆSX�oTڵ�=�o�x����k_Rp6��)��`r�!�~���@'��~@ '|�av�D^�Y/k�9�	;V��Ϲ�tZE�����u�+m�ݜ'gv|��a���'���x~83 ��.Hn8�E��~�\n͸�ta�ׇ5��#�i����R)�w��Sp�to�&���C���Հ\��c�k&���+��OȖ��~�ｄ�1~����� ;G0�c8Y�6�)�0�
2����I�8��u�N����"�Ĺ)��p6�V�ǄjV*�b>�ݻGGG�������s��#�̌�
w��H��*4�7����R�!?���m�X�	N>�$����:�2m����'��͆�3�/��MyP���
0�	�K.�E�Ӆ�L[�oc>��ׯO�T`
�?���� �q�K� -��!e���%N6�]Gee��Mar���� ??'�%�^����W0MI�H}3���p��X(M �5����	��E��H&8ubF>!��%�<�}����>� )�f�	`e��[i��1].�㹑/�c�֣-G���¤���ڢ� ���n[��D���ނ�a�_������X�� ���� � �d��=XZ����D��(y� �����ܹC@�o?|�cSό#�=���?a���ss�(�}n$9gm
%bM�Q<|�<������S�L��G��:�L�� 35�e���T�hL���c�[!��3�-0��_����TKs����a:���/^�6�����|������[����cSʜ�"2�B1���O��Gp��[�F�s��� 0��un�NS����J �ÁmM��D�~C��g�ѿDZ��n�9���%�U���#�\�|X�P�e�Qa�3޻C@���,p��ؖ���7�u �V��!�QK����K��+�߂��8��[X���&�J
�ZV!t)d(:�:Ёߑ1B�-;òo2N�	aI:;�c8QNn��	������r���O�o���a���kʸsvs��"�KL��'M�nY� �FP03��_߇�g'p�(�pw��ۊL����j�L'''��dr���G}b�$�VX�1��C�"� (eGfv0�y�k#�IW)æ��p��-�u�^�:��?=�ә3b�w����P<4�����$����҅�V
�,3���w`z�8� ���1\R��|��nߺM�~z���i)l�������f���\Թ\P�<��� �W?���qrx��Gpb�N1�i�G1�1���Wq�w?��7�miK[Z�� �l���i?�{����}�	��˯SE�A�I�n�h.���xj)���(��$M-��H��`�4����Oʧ'����m;�"��Y���1&�;����Ξ>���ǆ�4 �0����:ǎ��y~~^�T�vLG
A	K��<���g �4 ��z�+�-{���������X����#3i�2�� v?�5�y�k8]�|s`dΈ���{�& N�!߿G�~O���M�ܻ=���](_ig.W�(��5���ҝ$݆9��O;��:�_Mx�x4�g�"�Kff���W��U�+80�u���|��鷟_���{n݇���= 9��u����I��}�kr�������@��)���ԀA�{n�:�۷�Z����F-s���w��cYxZT	Aq� `���_ox�G�9���Wbi7A3�� ���у; �Cx����G0>|H&cg"�(�N�g���m��-]�����{>�n��u5 V�l@��6�]Ē-m�&2���������{_��__���O����!^���q��g�F��7�b��&Xl��g�F�y<wxpH`��ￇo���@I>����C����O�� ���L�QR����:䃐��
vv���O��}�����'�����!�z�)"S@`�1G�h8r~8uT&��C1SVt����}e�1�UA��9�ӷ�p~x�9�?��O��?�y
�퇰c���_�,F�ȧdԃ����}'�kMʬ�`�\�HN ?z�~���W?�Iv3�Gf�9?{/�OL;�έ�0??6�yF�q>��y]0R�۱IXC �}�B ����hg��w�87�k�}������+8����y���7X�OfvX���ۖ���ˡ�Ȗ���7"���;p�<�|�#����/�Sx���������_��0OlNe��:�+'d�~�f%�|n8��|A�;�"ay�$�yj=0�����o��z�ʖ;���n��/�������/ �s�F`#\��A��Y?d�kyjY������{8�s8���P>}	��X�6D���s��&0��S�Hӛ��̇4#�.�Q�0�j}9�����wH���?����[XQ��]�|���_�Wз�"ۅ�0���.��+љ���,k�T�S=z�����dӻp���������+����Y����� 7���G���8�Za_��E��.�5`�*F*��A�.�VX��Iؑ}f*4����ݧ0�?<;�'���"���m���X��&����_�wmiK[�Z�lE�=Ē�-�t}O_*x��Rd0����p~	��ë�Ó�!s8L��C8�ωI�.d.��q-�rX�rk��IgH�9G��pptHR���^>����B@Nw������ї�y�1��CPh���J:{�)��!]3����[p��+�=����{	/��FO��nAi`���2������s���"@�|��A���%���{��|qJ���м����s�������3(G�0/ǰ��o������~���kI�k_	e����2�&q6��5%��
�h3��� &����3���4��0����N�(�����߿G&��P�T��ѕ�"�Qԟ�H��
��Y�9gs�(��횾­[�)?�_z	/��[�B��	d��a1�EKd3i�Y�"Ӂ�����ϖ��E͵F� �E�</N.l���)	@�F�Y��Kt�g�<�F�4��l�X�K�"s��^4�NI�����@1�u��Q&�ŝ��W��x7���]���BD&�炛����]#�PǀVv�^�;d�W��	���>��A�/���O�����ŝ�%d%�&�+VѧX�,�+ʞn���u+.+�����u�Q�
k�N�0��ًW�l;��&�0a��Mv`�{�0I�~��ap�7�2_"K4��Q�[�z��>~����ش�.F��f=-��{�S�F9L�=���%<y�� �S���i�^��P�l��#M���܂@mC�;���|]���{`��l�!xW�gȽ)f�6�(�'O�3^�	Fd�`�������`����r�.�z 9jc`�GN���K��b!���7� �����_ôQ& ��+���4|����p��	����sx��)�)ӝ��G#�1����%�-��<�pzrNZ�Yg�Q6rY���Ch��Hط
*f37���h2���Cp|��Sx�&0��s}�[P�������G�2��N�+�����i�T���oK��x�\.U��1�d?7ݐ��c��-���ܥ<��j�iM�y
��J]���0��E�Հ\�h!���m�H�m�_��q�/�bfJ[�ȵ�%�j bx���a���u_�����`�`�{>������C--��qVcd�ΜoF�M�_�QX+T�`˲�����NO��30kt��� �w>�[_�G?�d���j
z)��,�� M�oH�9�����4M�&6p�0�{p������|����j���;"	��|fھ$�m�2�r�����ڕ�LMuFy+�lL���	<�
�˅A�� ����_`�� ػ+��Hj|d���$}�{s9/�^"I���.OJa�iv� �M_||~?�%�ߟ�� �4`|v���p���L�p��]�� �4N裈Z�M�v�'ӥ�<C�5~I�`���2��2@���cx����!�=�L�d�?�y�o�eH�ӟ��?i�����5Xn��N��~� �V��si��"B%�L�6G���7e��b���dK[z�$�����y`��dvhK�$����������+�
��,���3xq�n��3�01�O�#bj�̊��� ig^#UN�T�Ȥ��&�3O��+�%�(93�C��ܢ$I���ޅ�������wzz`���+����y���aqA��Z�ݲĆ`�w���?�� ���������ۻ��p��,��6� d��t�F����P�
3��s:�eM������W'prji�kh������������oAQF� NiƇ�*D���[�`�~�[���W砞�;��ffN�b	/_����4!諁��L�
�J�M��0����f>�O5���%X�������9��m���?���U~�3(�P�9�3el��X��h|�$n�5%��h��[y�E�$�\XH, �sd��� ) ���R+i
��f!�Xe�E۸�7�����;�31��.K�DZg��0��[Ó�@N����/�~~�<�K8� 2��)3L�x0�'a
�,�pa-
�o�4 �yF�Y))�A��� v@O��ѯ�����@�ڹ=����h�@�M���|7�v�w����.�x�´��=���|����g/`3�L$���!�\�v��FIR.�Gs�H0��V6� ~�0�t�>_�j�4}1qx�L=��� ���V�;�̌�;���}?��MgnghNU88�Ȁ�4 Z��܅�������v���:;����̱g�c�c��L�)ĵ�P0�%3*Kg6,av~J��1��b؜�f�n9؃����_���	��XaU�Y����	�VZ��r<�t���=X�+3-|�x��K!:��dw���>�t�� � ��\n��}�T�d��KǾe_2�:XF��n0X�Y�U�RH',�Km�t��/�ҎY�ˤ+�($�W�L��6���iD��Gp��]�|
��=x����_���cx=+`h�������S��tQ�L!�L���ґ!��M��)�ad�����/����#�@�c�]J��&C����fAs�l�oޒ�K�J�H�$�-�Y�A6ށ{��C��g���=8���`��[�K��`�Kd�,-a)�Z3+"寇6��|~N�Ѹ.0������Gf<<�(\��=�L� SR�r�%Z��-����E�5�`�}�ߴ���p�3�{�� N_���K��NNNaj@>�#�2��Q��T.j�����!��ϭ��T��O��f^M|��̳=X�E��1t�Ȫ�☲Qvy�����z+[�@��o�u��K޼��y�/y��FW%�K�-��Sq���j@>��~s� �!T�ߌ�~s&�֡���6ڐt�������D��l�$iuN?b~�g�`
�N������ɟ��w���`n�����b$0E�r4)��{�e"3��Z���z �[���/��_��>�;P�=�X�ͽ�؛�p��B@~��rK
{��/m�� ��9������������s�?����_���O@�d�xJ��ֹ^����5Vnԅ�hi����2���!�����=8+sX�~%j� �6W�eC�q[B��)p����|���2��|wtV�~����ٴ��\���PY����K:��0�@a�K\h��i�N�+G�������{0���}�{('�A�ކ��<-fN����\gUO΄ނ��O�߮����m{��6�g�U��_5��I���zMx$�+�J���ή�9�n�"�(������0���0=�����w��0�?��Wx��� ^����əwH+B	8FO�%iW@���a������߅۟�������%;��P��<Z�ct�3�A�ٞ�����2�\�[���:,�<����L#z�x������7�^�d��J�G㡴� �܄3��9���-ܾ���p��W��߇��XvI��D���Ȥ��nΡ\��^lx���_��ٙ{?a�u0�q���� �x�ʳ�p��w�쇿�~����b�K�9h�Đ���mVْ��y95Q���_���Gp��s|N�(�]���	dEyF24���Pk@�u��Z�j��[�Bo����enK��6x��#ե:/q3'��\"т\9����t䍟@��h�]<
�u�1�Zzo6��)���!F�Qk�|����ډ�ɜΑ������|����Jî�`��[p{�!|�+X>�f�ë�/A/W W��B(B�*Hc�H׃�)c �<2|��u�cS��a�9fa��Fd���Xy2�����������E�c���<&ѮM63��P�s���LMa8���Cx��7�ѯ�����������A��t��G�F�z�9=�ľ"�q��2��DL͵v܏G;,�)�D����'�Aa���3��ْ�V &x�0�����djF�a��g��<f@������4��� >��{����G�����2��h�b gf��lό��a����ƗL,]�N�h�:����E��?]�|��'PsȯiХ�f�^���FQ��\P�u/�E����o������Ɉ�n@&��!h�{��ܺ�������Y��S��C�K?G��!(���Tĩl��>%8ҳn#��$WL��������$�qƕ�C�*2���F�I�_$Hq���fg����_�]Ԩ�_��v����Z�7+�4�o�B��af�<)����a|@L���G��A�����0���s�M�e�x���.�5��xߔ=�e64�2Q+�6��i��Y�1��(̜�ĸe*�s�1D�I���U������E7a��濰�O糵5g��")z�BFf��^�#e=�aޢҀ�s��4�Y9yt����/N�`u��vM{h�|E������o�cJYC��h��6h���B0�[!js#A��(���gJ.W{�t���}� 4��&��X}ϜnJ��E�>7 d�&PS3�1̭�1����O!����|�N�Bq�Q�N(��� D�񲻻�����;00@~��3��^!lD;��0�π�B���ru�lz�L�3�'�7WoLW�5U���O	ɤ�h��I��O���z�r<M��6���6�o��*��I5࠶Ҫ���v�k_��V3w�U�+�3�̈��.�pҺ5����w9���R>�~�u骣jm5  ��D�+��LpՔ��M^�����R�g�=�v@������v�tK�o��Dy��GkM�5>;��=�ȟ\��UK�Ȯ@f*��\��uc 9�E[;~��/j@(��abI<"��*M|�&��i���.$a����M���_\56�R����'7쟆O��	ѿqt�A�%ޚ�A��!�_��OX0 �����W��U��K�2��*����ֱy�\��i���Qs1p���$I�m�lH+�^�G`F�0���M�~����D,�E�tv�o���ʏ0Ђ0`$�?4�㲞�
�?38�����o�"&�ľ�L����s^
���%���$'�\�U �`,v�/�{_i�~%���;�һ�ʋ�i�����r�ˡRiO���"���
N����{X�<�_�z)$�:m�%SY�@P�WR��4��3�Y⁜�@��Ch����T�F���������QT	}�!W�@8���ů[/Ȏ��ڛ��s�r����F�@3�>�ȌL�&�r��x!
x���_�|�&�� $sO�l�w���*��h>�6�J2���?������i��c�wS����?%cԵ��Q(]eO�ϡ�f�@�aV4��Ɣ�e��~ {{�^��Ն�� J�C��G@�ד-Rq݈�&		3Hx�f�����-��ry����ȋ<��ÃӋ�'0S+
�+���i5�%i�%Ey�P'�T��,��/$�d�h[�ڮ9"�cpߧn��-�m9�Kյ��k��=��
�@x��\���M������\���o����K`�H�&����M_����6� s1ֽ���� ��S;�)=�����G1*j�I��<���s)j��'٩liufcNI��NJK~�ɲJ�\:����5"[.!�L��cb;1�F���N���n&&xߛ�e�I_b�	}u&����WN��ц��BjA���X����J^��2s�	:��˅&�q$�3�ٰQ�Y�O^-m45�l	��YTe��d37�����t�޷I�z����� ��@-�bT�o^�dJP�w������h���m&R���2>�"�'�zQ�z|r���y�lq�z-�p7p���]���7�^ r�_~Bm2F������#�ކ509ba��j1�YP��::�mأ���2�|�g!�6�6ZYw-r�`F���(���J��BR�0�����KG&2W)���O��7�Mm��(����b�xĸgU�t�nD-G��aV%��
ծ)���s�b�P�_Yk98�V}Ύ�-cX�?K�6�O/�g��ٚ�#(<ՙ���MCd�f�
�b� s������H��p8�_j굶��k5W��������]�)�b���A]ؿM
�Ŧ�_S׫K�C�ǽ̳P�Dm�k*�Yb����Cl���{�@�G
���7f�ܬ������{�m�c�OHh`�6��]B}.�I��}���/n���?������
�t���߅v9A��b�G8M�{i���_�>ʅ�F˛T�o�I�sQ��ՀlH��%;"��Ro�030�Cg�U�����S���I(��'��ǜlHR����(�&ᤢ"��ӵ�p���N&=�������]�so,��ѱ����Ë�A�2#)�޿�����' �ZelB���˷�*:k�C'���'�#��ot�:"�G�у��w�1S@�_��I���qd�Z�12l�X1LA��V��=3Ir��l���_\I�e�5]$ާ~k'-&XW,=>8��F��������x|\<������ �
O�C��>mȆTgAgdL��Y��b�J��0(�C2MX&ʻt�Fy!�	�I	 �/�䬕�DbM���碱@��H����������rh'����rf:���#��99�:Pz��mc�׽r��q�C��bw39k18��ō~1���V��/�~TTfʅe�LK�5�I�M��"�n���M��ZvI�z�#kz.Կ׋*��;LG4z Cx��3������W�Lm�̕2��y��0�w���2�]�2ҿ^��v!(qo_���(�Z�&ig��b�|U��̮ٞ��۠ ���~�DfX��2� ��� $gn����;���iCx���s+��ps�h2���j����c�������!!ʯ%6Z��*�w)b)滍�[.w��1��f��$ !:ϵ����->�қ �>�����|���#�C��`vJ�zD��6�iW�m�n͟���|�RR��>m��I�������S�����;��`�������|߄��z�r���6�p D��%���6N���G
.{n��f�??.���9mG��kQ����� �m�,^�t�����M���O����'�(oS������Ԧ�
��ҁ �w�����V8?zYXJ�́���@����?&kC�m4:�k<͡`�_�H���3ؽ $���]QfC�@a|��C��˭C)�LX�5����2�s��o�´R+X	S=�r��}3����03��,0d�pT�[Z��F=����S��V��c�!� �����|����9�G��ځ8:_I�d�$v��^-���ljM��_duLt�TyL�5s�0}U��}�:��oIb��0��2�SE��{��!5[��:	 ͞n;�}�B��ZG^P^ĥve~��Z����*�}�6�ܘu��m�1��J����>8K �������Qܨ�����;�s����ͳ���V�b7k�cI��3�\�fH�ڍ܂�zs��tk�GaY��}0��vm���\��0�6�A�m/�׾o�z����$z��r�o�e�F��h|�}/�4�j���[����!ݯ�� 3.���+Im�@�U`���3up�g�d$$���lt���SjI^�'��! iY�D���`���ۢ! Z��=�����3�;�o5.�.Q�o�W�5�-��/Ԩ͹�bpA���S��},ǥ搫!.Z�y����NP̂f��X���5ǒ��#��q]5)�j@"��y��VY���ρ�1��#�blX#ʞ���l�f�f��B���^��s�yt8�1��`�#�K�����oѪL���θ�9RN�/CYM�2��p�U�1ɊaN$��U�Yf̸'�2^�#����@��9����tb���om�Ӹ̎)�1���_c��̙O*`l���z����N�M4�K�(���F���~��dj�lO���u�Mz�>���+���,I�VP�*hw�gκ���#.�f��}�����(	�����5��`��J㤼Ǖ��(㲼WC�̠��|������0b�D�Ɣ�q�����U3��r]@�#!=�q)��0�>sN�o�0��[��i)�����L�����O��D�͏������c<G�u���4�9nӄ$v���L��Q���acB����p��nG̳�T#�qL�e?�;oi-�Fd���+�}����&�l��W˨j���u<�nw	���f��#����Mؽ47㬄����Rb���Z��
�∈���kw7�=�'|��3U�����a���v2��0++FQR�+�Ϡ4�X1�ӧ �%���
�2��hh�2w�l]3Yf���7��s�e%wŌP�?�[��- ��D�/]�g���v�l��y�u���x�H#䤦X�5U¯/3t���ޠ��� ;@Ŀ��M˚�Tad}�tIŢ�2߲�=oؔ��S]�҈��Fr�Ը*Î;NU�h|u|�_�7�x#���Q?#��3ٛPJ�0Q�� �cZvE�k�+C_զ�5�u�jE�!���)! ���y��R=*��\�`ʬ��+aD?�ujh|���ލ���q���=� ��5��� #>����}S�B
G����
�X��zFA��)ZvG]j,���D���zT��q�s]����� 8IT�R�}�E�!^C6�jf�ycS���W�6ޯ�}�#h�΅����b��EL�J���l{�/0P�ڑ�;:����j�}�;h�|����� �P�` �f-86��̓raޯ�k%֣��J;D���D����b�����D�@��Ւ�KB���f��(f0;��^|��,�X����c�D\�A:��aZ�s%X�.>>�r��T�PC�r�b㭰�l�@�&1��:v�o�L�7�?���Pu-���*Q+YT��V#�}��
7믐{R�Xl�2'=	_�cТ���N]@҂Y��wdr��>C��`w<��������^�R��^��d5d8�W�T��k���2���o3�f{�&fm�����93`U�&l]��g>���+�Ick��f�=; �{Mm5-�l������oP!�h>?ր��&F��x�k��aDU�f�=�+5^��B5��Gl�N�x�]�Ի��Ԝ������~�U���/�6,�>l��mp[�^��,�o�{�^#��싆��f{���f@�`8�QV����O 3<�(O�8�@�߲*}묰SS.(��z��:c�?�i]d�{]���r�< ע�)B�ܘ�\i�ZU�XJE��$؁�K�T��Pݥ�̅V�%�N�`<����0sx��@�_B�Ma>���0�N`������a������c�p���m.n�DJ��.��en'�ْc&\��4��U�"��D*�BlR毇��.i��B�)��\T�vG��n|�"��0��t�6g����]k�(n��	�1��l����� ���=�U:f92��0�C\ՠ:Ni��&�=0���+[��Nj'��u�4_U��24=���鍡ݴ�>��
��X��G5nt����m��a��`��3]K���.Y�1�l0`
Rㅶ�6 �Bq{�V5��k^�r������)���g��kŸ���+׭ʤ2�@��VpJg����o����L�B��>�5�^s����P��n@�폛�մ���9u�i`hr��z��W�ȻV�����}&�"�7��FS�)����3k�m�ScE "�4<�c>52�3k �w�����z*ݜ�x��0���/0��?W��>�2���I�a��[�'�lRyX_P�'a�оjށ��ab���0��6�M�sG�?�r�����������Y��.˲��v��"��y���v�; �y��Bv���*��,�p�ҀT�����c�s�
�i�f��$���2��|e�wqB�ܹ���{^,`nЖ��t�}V �[�,��S8[c{ ;I D�
`89��}���~�g�!T���?#4a*Z��x�����&Y�Q�b�>=�;3T����T��X��:�RXg^�2���_�c�"���l��^��f�F����jJ�769b}��A�[o4Rd���꽲c=^(y��<1<l���&QcL);���$*  ���ub3 �1�|sOr_9ئ�LG����1�`��D�|�SZB(�����)�"���v>u�m��wmb�dM���U^��p}��C��t0�t��&V�?5^��7~R5�v��8f�2Y�̆�Ĉuh,Q�����.�`M�C@���U������) �<(����u��:�j�k�
��ʉ��v��fr�$���e���.eQ&��Y�_�� �@z���Or�'Q������E/��~��G�z�A(��H�V�aߊ����z��c��$�9�$�T��(eA0PR�
�Mӹ*�$��<�/���^Ts$�|z}�.;���������ʥ/PÀY�_����{Z�7Ӏ��w�	�$�T�XeG��R�a�M#8t�^��СJ_����h
ӡ0H�U�L�r��e�vAg%�����9��Mj)ˠj�VIZ*�� b� ��z��oO��4��u�SQ{aT��/`tS�=��WT���k����������c ����mDc�If2%�NP*�7A���>�ޑlBc�h>�@��q���/K���wB%:���82�na������W�Q������GR�Pt΋zAW՚@~%*�{N�ԀD]u�7�|X=/�F�����y�<[����T�f���A�5���u�z����J��HE=m^�4��G�E똠����W��V"����U>���Z:]z�����'bN���>��;�M�� M,A'�����W�I8u�	��Wi�T{���xeWk_p֮��1W'���S�s+���n�������u,�
�5��	��GÄX7�w�q������Y;�X�V��n����ң������|W=����l�	�����"���������ѰQ'>���P��Ln��!
�TF���V�7*L%��	�_��FyD�H0-���tI�m���*"��C@�I��"�@���.�@�w���ga����r�5� ����wD>�X,�:X�6�������g�����B
	X���=�/�i����xK��/N φ���؅�jk�prP�6Wx���w*I2_��2�1ڕ	�e"PIV���|ePe5(���X�CS��u�=��s[��Z�T�E��rj�F�����Ty��f��P�v��t(��EZ6�|M �
L����KФ�v&1X	��g�`����C��V�&*�X�G���
ة�	X�W��`��F�*F�����kh��V����Ac�ה�=eb՘�����7��k�h����=?�L$��5�&�5W�iM���`��$���o=,��x�v�|4}&l��.W[�k5eCSҶNUN�q��Wƌ�W�(Nt�s�pV>vM@E+���G���m��F&Xi�Ϧ&X�h��׷E� �l�p����:%��SQ���n0��r�n�W�Q�Qc�L;~/[MX�h<�`]`���n�ui��W����8�Μ)��B�π�M�sS���0� ��E ؤ�����~Z#��n6�U��r�#�<h��<'��<,�g�.��k�\!u>��dY��Nqi#4�h����`����S�Ďe������O$��˝L&Bdԉ�5?acѓ���ݷ�T����t�)�����f/_�E� �r��E�6��I"��r���3ݦ��u������s�T1�I�dX^�M�����Z���ME��UN:\[	�U%���� ��ҁ���o:��7�P�C�����3�l�VIaU(я�m��$��Ԓi\�Ȟ�)��U������2bH@c�uΌz�te����_�ɉ�:0��ʯ�n٭3�.  ��3qh�T� |*_�F��d�b�zB�.�ͤ�������c@Zi���$\5"	uU��TZ�@��E]v���rM��|D�o��f؍EQ
h�+�ѓZ.���&W��fz��A=Nb-�����,+@�L����6U�V�Pc%�0����'z[L}N�U���G��;��͛U��}�4���4�=`��o�_ƻ>���BM*������Z�(�K����F��h��'��D����0�m��},P(����+�r���C�g��)Ȯ�_OB�-/�Q9PHV�K�*���Gh�B�Zذ ��Jۍ�±�e��6��eQ�x.�|��p1�� ��ʫW�`<���t���<���0�r>�B�v���i@|������?љ������@�����N��)"zd������$5���NϞ�P��Mf	�e6ܥ�UF�IlŪ��J�V��t�ʜ�bX�va_C��*�/�(4�:���'���2�l�4��U_"�Ku���a=Dc	O-1��W��Ss1xa��pRkgn�x# �&�-|}����#W]����#y�@V��-��Ϊq_r�����
�v����w?�J<�9�f�pw��ni�T��M�cЧ�ɱ�I��A��۔zgi�X\?f���9�Uݧ�Q�(J^u{l"�^�R1С#xt��=�,R�b(: ����2�߫� �k;|��y��=��Ao��Q�n\gK�d�58�Toޣ�0�zOO�J�}4��:V�ܢ�z&Vd*��%���tu_y1�b��/���؇02;]��	����%ޱ����<�敧��U����ly�\��u4�������`Uψ�ܻ��ӡ�<-�>�J"�a���;���Q�wTK7���e�s�G�t뗷�Ѥb� ���V�2�) n�P�5�3�<1�L�_?wvv��wD��µ�a0� �'~�O�sc���83ze��9� ����3�*0���Q��/�3{���K��hi�q��FtF?�,%���QV/�x���S����D�px�6ٜM �ր��x@D#�T�ҏջ�.��!u?Gk�5'�7CYr�H%�4�s���|j���A��MM僙?�����;�	='`����i]�E�u��&RjC�t	c���:�K�������>�(O  ���QtK�����vj��	�&�MpR�]G/�L;U���IU�L��.�-vd&[n�${^hײ�ǳ�~�n����W�iR����>nh������̼GUP2d 7K����;R�JQ�D�;�-�&�5ҳ�/���t9���5��A5�"F,��ϭ�&/���oj��=5cA�N�DUy�x�M,z�����Z��"2tT�Q��Cv/�TϏGx�<����v�ש�^]��*�T�Voٱ^֤�0<�z�*y8A����UL����?�N�M�!@w�ae޾(/�\9a���iO����ra}���޽�5�!�`k�������2��<�[4�Z�� ����|s+�m��D���;G��0��28</�r��X�o�U�l�K��OQ<�$
�g�mԐa<�Bf@H��58�c Rm&�b����N ����J�ژ� ��\�-��"��~o�`o�	.r�.�az�}��ZcU� u}���_�!�<����F[�)o�]feOK�䆫K��r��I�Һ! ���e��֫cq�7<�QkcV����oӆ��l�cJI��gK�M:��h�nM �b�������%���PK�A�F�&@�F����U�=��}�RN��S`����N��yĶ��t8��ڇpސ��Rd���G�|��ïÌX>�˦L�L����	$Z	�v mNS
�����^�5����셁?���c���^P��j$��OSl�\?=߲?��e���I[lA��t�t��BWV'Z�/Zbv��ϼ���J�d����a�<�|d
�p~zl�,>��T�ù�
�s>!p���(��Ѩq�
��]��8�O�;�u�d÷BQW��a��9�Ⱦ)n`T1!��3
�����;�����u�6骑$]�;:��rŀ��}���,�D��hc6C��&sI�ͳ3W�N�f��/x��m*@���E��_����1m_��v�Ou�Qm�P����N��)b:|��X�l�~t�
����ˣ1������WmNQr�.b;y�b���%v- 
�Sׇ��b�}	ڲ�~��vK�ڜ�����o��C@��q�XC�.�		rw�z��Y��?m�����we$1�� #ߠ���+%�h�k]� �'�P��4u�e��&��QY2��E&5��-~L}Q�ڨs\��^�O�繘n�냪���]�N�K!j�:	A�����	���Qh�Mϧ�&_1��+v2o^�� ��ɣ��j���6����� 1�����Ws���X��ck���l
�5s�p�u(���S�y���z�E)��Uӵр���84�Oq������N����A���?q _�� �������ŵ�]`�/�q�M�
�J�M?IhKT�_[Ie��UR�F
 +)�O��Bt{���FY�m��)�16��R�8n69�5��\Cr��ͼ;JF+E�n���@����vT��@�i��ןd�K��^���j\ǏZ��uQ��J���܎�U�K�K����Y�e�ק:�<w-����i<�s=��� N;�[��`I�� ����4�<+�\���Y��3G��BlE?Een�*hoL����<�l���Z���kB�?�7��4�+���������m�樫�8���[�0e-A��T�����iR��＿�ſ�-�4��w�k���: i1�eQS�Ѥ8�L�|�x����=h�`MU�:7-`Ȱ�	����Q��q�^���NXx�u�+���;����}��u��wE����}=�Q�4.m�Zb�%�|o0������e����l:XU���MbG�di�	�O��Ν]m�j��T�e�V@�m?�	�'�AF�'4� Ν'#IL'?�s*�&X1Qt	n�M��h_�Q�j�&0��+�Hmr��:��wkXg�	��t���:� 8��/WFIҿ��N�筣��:S߶9z}2���q�z@)���W����w)��f�O��~.�������m��X&6�J�ӥ1��tV�aE3�S��vo�y.e�Hz_�8��-f�׏^�V]�1���6S�|0:�y�J��t�d6/��q�m���Y��E���gR����(�)��C����	��&F"�������r}$Ds�JF�ka@���l��q��%�fXgj������>TCV����;��h���9�~d��h�>�����z�B���5����. ��׾�w�Z��MI �{�O��y����<��X O���.��BT����f�灃���Gd��S�Iһ6�z� �ox��`ӫ6 /�m��'���<!:X��w�}�ʌ�$H��� ̈́�C/�V�$�viJ�� �l����b��h3i5+( �?
3Q][i�	��NM�썀G���ԣ��I$"ߙ�9��x��9���WTI��Y�f�T QSk$��k�(WK�0Eaø�h�_��byI"+��xC���gI��=o���3�΃A��7&ތ�1WlM���qo��1T\j-�jJ�j���HI��w��� J���FL�;U�`x�=�0T�X��S5b�Q�IH�"�1���!"�)��C��8o	�3�/=�ՙx\Q�~J����>�������n����������☔)��=G0?m�f�a=�y�*�gL�P�{^/�i���
�Ȝ��a�o�盘�B�g�Ǉe���*�Z�xɪ�Z?���b@i�*�}H+��?�֐ꇫ3Y#�=}ݽ܍�Hx��\�<=��w����D{NO�6�Y�hV���V����Ԛ[�j'x��`��)H̛njbu�hc rա�|�͡|jC�}�hn�G���>vww�����_��V�X9�y�Am6s_� ='+k��aL)ʆ�A�"#g��dK�j7�(�.�V��#��c�E(�u/�R)B�`��0�Xl:�e���;�.�&J�~�D����e�2��_�z���!� P�� ����Mё�N5��XB�w�^�j�&x���kR*���Ɣ!@�l+��޵m�d0C[`��ǅ0��3/=Qv��y��*�\m���mqj��<���D{��q�G���h�(�J0l:q>~^c�2��UO����#��L_hB�\��"�gXW7�j	q�	�o�j�̚Z*��Ք�m��pb��hleQ{64JQͫ�q��V	�<�]�	��Y�F�����>��_��/`�ۖ��c_hX@��6��ĞA�⹖�25m��G��FM�� (�o�(v	�YJ��c������ڸ}:�g��G-	���D��m:]�j5�h߿{�᪺>'�Z�µ��{�����*�wTN��/&�Q"-,
�?����x�x|��+���l����1]���;׀�(n�8J@LmRe��e��O,�Ϟ��c�C�ցbI'x��U�6�ڂ�ϖ��Eű�z6h�~U{Zs �I�	�p�&^�ty)z��4U��.(����ΠJH��� ���/�n��ƥCB,�2�ƙ�D�-%�>�Ukf׸���SA��&�'�B�~C����y2���=��Я�����>-	�Ƅ*%�q}@I���~��4�{�m����aS��������Jj{J�$���FQz*&�]S �o����%T�˴l�uL�A���P�CW�I�����W��t<�g)p�~�i��T���R�^F6 H2�o�� �Q��2@6��=��G#��U��x����'%�j���j�°&��7���R*M�.�!��Fb�u5�d���Rjc�O�����^�R�oZ�U�: �XT�&�&߬��???'��L;��N@�����o ͧ�P)�t)���Wy�B�b]?k+ �!���T_��H˲) ImP�B&���4�����p��N�6��1�Y��f��H"�o&H1�<j�`��-zj<�t���"<��0`���o�-1��P.
@R&��20S�?�>��`������ְ8쥤OEd��n�,��SP�H�g��.�{m����ˉ��|� kJ�c�w ��$���Om�`�( Ybo�}HFZK�_�`��1��� d�奂��4�K���L�7]/6^�.��H �>_�������H�P��I�bHm�'j@����O���Ӻ ���E!w2����Ik�pʉ%����I��V_Ai�Xu�n&�^P~�A� ʑ)z��$E�wk,`I �PV����G�&lD��E[�80�OEJ���l�z�1z�1���`�L���7Ș��l���@h7>��T�J�~hr�*Z��>~خ�KHl��.��20��X��?1`�ˋ5YC#m�	�� �:�/)�u֟ @t�?���z��5j`��� �WA�?�M&��D�:l��\s��G��c'�"�w}���2d�� $��*������[��3����Q�0)i�}�7�l�~1@�(�F��'#^�O�<�*�l&�m �T�x���w��>5� �S9��'�Xh�y=�e��������HQ�����P�� ~��x� I|?;����^�5 ��d�7H�Ym�A�M�Ɔ�u�M��:��M�yX;�&�hZ!G��q�������D pD(����fe���O�2�=&X.`�>���N��L�}��^�y�>m���a����Pڜ*���>W�Ӧ�@$�Y-�}�K`ml��7Ll�B�����		k(DĀ������_�yڟ��D�!1��(]\_��{[Teʠ�3Ѫo���Ϙd�c�hϘR&�A����}SȠ�����ZJJ������v<��_hbx7
�H�Q����s�D(Z`�,�ktB`�j�F^��3% ���հ�6�_��(����*7�o[ ��g����~�m��F�w~G�pm��N������FQ,xStG:��>}%jH\���|���#C������g�!��W���!zwv�M	vjCtN}�K�Ø8�13)�#����p��ҡML(9t��ǁÜ�\S���Z��r�'�Amf�������9��\Ƞ��9����uy{I���4!IDz���"'u?TQ��b��	Vy���xP����rY�C��-�Ar�g#���Zb}�6c���e��<�� ��Û����E��Tb�zY҃�# R�A@��Ӻ �W��z$h,i�Q�!$��XF�1Y�o�����ۇ�~N_��-�7��XB�"A迟�/�	�#��o��O��q�7��M�JR#6�)�� S��l� y&'Ү�Go��t剹6�q�Mo|��]��Ć1�||R��E���;�� `�g�l;Ǿ6(���5�}�\4$������)����N��ٿI��"t�E������́Cv	!ܻ�lo�>)�{3H\)]���	��u��OM�����$����(��q|� d]�z�>e��T՛%�3�A'l֙o����X��������hD��7q���5mfX3�)�/����y���f�@¾�YЅH\���Z�d	=m|Q&,��'M�H�?EQ���nS rQ���Z���&��5�0�6�f�t�+ �5�-U�	'�����4�S���p�+@Z���M5`���4<oq5}��O��������c�d2z#JWh�)�.�(�����&�O	(����w��<6N���j�N���Xw��<�ǖ|� o[=����E��q�9�Y2�~�?6�ByN˪�-�b��o\�t�$E�=zN�>Y�;�6(�'C6l.i��ܶĹ��1a����I��8�[��������03�` � !z�����Z�n��������?��xbPR�{��H�EI%�~������i�]��o~yn֜�S�U�U��~�FO����c�;�e��w�1]_\P�p��irA�u}6D�~��8��������C�bM�Zk���EcA�^4{������6d���T{��"�5c4j�pcY���vM�W���`�6x������
��-��4`�[Ś���7U�brw��j�-�i���\��2`+�'M���]��kP� �w�������ͻz$J^����1)��0	�,U�|����V�p���Ug������z��*��}�k��u�5>靟Kk#������k�w�@�e̯&$��k���թ$��C�B�
���A(���E�Xs�sC'*wf�c��l�޹��>YӃ|�G��񅀬1?��jT޸5���I+dh��G=�u��������5��6n�H]�Q�� !>|(���q�2�N�fݖ4��.,-h�mf�����A�H>��i1�[��v���Ɔ��&�^cu-�{>j�| ���+�WF���۽Knk�k��a;z?�z	Ȯ�w��n ���.���\�[������]u�q��G��l���i�*\�V�a��$�G��I@��.�^
��A�ƅ��\pQj���SލJ�[�5��Z;��w��nE�%!�w� 	���܊��Z��DW�VI�c{����+���o7�K���Il���K��$7;}o�������9�s�e�]jk��J܍�W5+eװY��� Ai�������Ͷ�*�*��]i����H�6t-��ϯ^��^[[vUܒ��v��N�(	�y�w�|lU @�L$�ID����f[}�f��V`��JCf�_5��:;���l�$��V�I�[_�����kLA���}�E^����Z=�n��uH�fa=d�'!�>	�U�P&�
�d��,�%�k%��\8i�C�t�����Q�����,#������}=�K�^�k�ж��Z�S�����sn��i��1�j�%�޸��Ñ����][aS	Hk�F�����7������%������]}����e4<�ާ��jy�ؤ�(�j���m�(լ[��U��j_��=t^��U�V�a�����Ç��{�Ԁ�t�	50g����P�>�>|����ǎ�n�!>|4��nW��O@|���Ç;>��a�_g�xB�v�-G@Z��u���i.e�3�
.�f�V4{|����j��o�:��t��	�j��8[[�[�}g{��ۭQ�n1 톭S���7�Fc4�����:�/�ъ����ɩ57+?�c��c?�/�A>��~h�>�V{R`sky%l9�Ç>|��ᣵ��X������Ç>|��$d� �ͳt�" �Xч>|���c��g���X����]��E�|^ϡz�Fr�z�ֺ�V3ڵ4�����^��w��n�j�Z��h��F��j�F۳���=��=j�_�x�b����ըў��{��b�Z�)�՟�=����l�����6�����8�J�cHK��J@�*���gUs���4���?�X�xi�;vL�z��6�E��c�����M�m�vF��9v��`��u;՞���b�4��y�} [-(���🗏�{��^�o}m7�?͎׍ �%��2���L�ވ�ŰQ��
��h1�������Æ��k�Oͺ솹�Y<m�+��OB��j�zg��' [��p>��a���e���Qjy@��ӛ�]�[;�J7r~�I�����`|؄d'b�	��S��Mi*iL7ӽ�l�C�u��9h��^TZ�lp���z�ڮZ�1�扯���=����za�K�:3k���1W�9oE�{�+͏vug[ڲ���w�͑�$���#�Hٸ�cU�~W#,��1h�F5��̀�5?h-'<�/��=&5������#����q�9ụ���[�@o4���kń�:~��Y�	K�1J��+y�*��dm�I��B���K>��le�M�1�-*a�	�����۽��t�5��yj�X68f�@7�O��X��c�m�����h�𞯖`��4ǫT��68|oN�Юy�c�A0�<��4e��r�g�ה��c���}�4�4C>v���Sɗ?��|C�Qy�RwԽ�V�8��7�`��Yg*��M>l�7K`���������f2�Uv���^?O�hW�hW����H$�} �D�V�ݧ��F���c��p7����	�.���ox	@���m�h�&�8��a�Py�-yY�z�1T&SIR��e%�s^YY)_��'[�_��|Y�a��v�\�?�&�I!��XLȅn>�} �%��$�>v7��;�| M���@���V{��m�J׻�17Zo/���4n�Lw�,֪�l�L���j�a�A`K�T���U.SM�o��x߷_�g�^6Cú��'ݹ*y��������j.�E��~ގ���c;�C?��FkF��mO��V���hw��FϧvP��N�Re#_�ho{<�";���� ��:;;�^2��/���v���6č�k��/�CQ+�F�͢���+�jwLO��og��Wk���D��IA�{@|l(gg�f�A3����VB~@o���4����ga<������>������g��J�p-����q�(�	�������~%�WQ5J��ZFr=��n����n���)�U��Pr�$T�K	��U��	�z���nu�t�۩�B����P�@�5agjtWRGmτ����6�=���Yz	����m�h6���X�w�kt��*Գ`�V;˖~_	H%�N����e�s(�х��%��`��=�o{l7�Qxcn�%���
�<O�_zbC	��|OI��)�����XlVּ��?�I�N$!>��5�kC���;�J��k�|�_%kIb���$�	Q�����]���SI�Wk�ٱ�<Z��WOZ\oV.�Ok_�x�F�ހz;ݰ�v�q�nh,5��D�������t7nN����b����SP����;<9u�F5�ݐ��ؾ5������f�fǘ4��7�#��v����~��m5���W+�_Nm{=.v�a�8y��Tx�j�����o�l�iX�Ojivk�q���i�<ܻ>5��T����m�g�����3�����Z�`��v��է+�k��ˍ������cU��_��+��1z,����Je|6)��H�� VE���q����}�y�R�F����>7[�YÔ=�c-��g��Fퟕb�6�=Pi�]��j)*���H����>O���^|�N�{@|��E��TL0Lt��ޱ�]I�8�F��f�Ѡ���W��iÞ<�-���۩�A�`{4k��ڻ����Z��z\��i6kP5[	x�t�B��jcЖP����?  6��Y��4�Y�h�Hư�a��f��>��cA3\�D�δ�dڻ� &xߖc�mԐU��,�� v �7����M��U�<�������VF�F�{��KԳ���,�a���G��y%Y뽗z3-��PO��B�F^+����H�ć�]{��cAl�W���j$��5X������4����Zݱ�-^[�e������#y�eP�P+���hV�UK��۠��|U�	��ՠ߷�;��;�h=F�7�A�d�������1�m+��z��M�k��_����h6�d!�bt��j�z=�mt�uUM�݂��h���	^�4����F{%�f&�5�^ԣ���ة0q,͠d�1z�:.�u�A�9|�R��7�%(*��~��>���J��**��J5U��4���-߳]?Ǝm�4����Q8��Q����}V"D8�-��ez���U��٨��^^	���>j�AT�s����^� ���Ưz��xvl��#|�~>v��Z�ܻ��}R����h@7#���<!������ �=�ytnk��s�}/�{_��t6{�F������kv��C����H�J=�5v��<��z����+�T��J<�ּ��{@j58nZw�ڝ�����F�������t1�	�ZA����k��6uR����B�x�x �tG��֥�	]</����0�5;ȭ���_��������5� ;�[�r���%t��%f��W����~��Ɏ��W���t���?�:�<x�R%�}��EG�~����hǊ�h[�Tb~�Mo�+����8��h�Ƶ��� �G���vq��~Gb�z>^�η:V�m$Ղ׮�6~�N@j���k�^h�	2�^��R�7�.e�P Ɲw�ԖJ�Aa���D����T�N:�<z�ji|ׂ=��0E%��V�W��Ə����z����B;����`�Yj�`^o�����ٙ��:^�Yk� ���ݠ�W�h��w�^?�c�R&�F=�����@�q���&:v?��Y�Ju�R�S�{��A���7������L> ;����똴����΂���Mm!ֺ`�$Rz꿷���?�h�
�y��ͦ��lT�2�ά�F�����AT�Lxw>���-oXώ�Z�G��*�����i�?�G�pؤB�:�ڰ�JY��P�g��$���?�! k�g{�*Ցi6+�M�#�4��o {�o��Ba�7�!!�YQrQ�k�5�u��޿z�o�@��8jv��>g�}�\�f�x7��B���:������o.o:�y�v	��:g�[���[���W�U�Y\=^-M�� �bf=�7��f"�M�z��o�]J�}�Z_�68�ϭ�o��B�ƙN*���Sǡ^�G&�6o&�Mz3d���tGT�x���n�jƆ��o�� �2�F{�ߕ
	�3���%4�<��������x��g-/H�_z�K�_�T���5m�g��|�}^�<�7P�A���
�z�lYD��F������}���h�x\uE���nf�}Pϣ�������9E艹�y����Պ�TQ�M�9��1��=�+�;�&X��W=ϣ����]�gm�ӛ����ݞ+�>�u�O������YW'95xp���4 M'r4�z�4� ��`�;�ؚ��z�8W���;*�Q����\�ී0 j��o-,�ש��5�:���bc-��z�~�,p�"��Tj�J��&0�[kL](�~[v���P-���ߵ���w���n����7�7c{J�~+�5+]���g�7%J^rc�����sN=�ǃ޿*(��J�㬶C�=�
����=���RJu�:��AZz~j14��Nv�.��lug��VSVχ.5h=;SE�|��BP���Cw���x��ǡ��TkB�z`�^�s���Nt�4K߯u|oa�J�~N��*y4mؓ�v0 ��Z�|��U��P�D�s�MV�#��K(j=�J�0�8��ഽ��64l��m@x�ю�Z�qc�}틺�h_�^���:��׳���9��>^��������,�!��l'"i�9�dg��7��;���= v�G ��K-�`	�.�����q�"�������;x� ��cE=���h�٨4�k-��v�1��0nUe꭬&ͱ%A��g�Vk�FQm|����̫�Ux�R�R�Gw�m�M�`��6?6#�m�J�#;���~��nl��?[re{J��TJ�`Kx7��?X�!�T�FWW�|NI���J��z`gH������������I}����O�#U��TJ.}c�m��Y)��H$��m��{��/�u�q�rK�;��z�����?N�N�����]�~]~�?��������|ե��Գ��.��5t��~�]Ƶ���c>6���j*��{�=��Z�Z;߿z0�V�aȖ-�F�w��ҳV��=I�3��E��Øl6&�6z���=IՎ�� b@���v �]������Z�z�T��(�j(��)v/�\��y;��Z�Z݇�Y?��~��e?�J^o�8�V w���A�*��܂���P���J��%UX��o��*]o��Uu�߳m�f�f�����1]i�n������|T������N����/�۷�������a�2��;����O�g�x�\Œ���^LMڠ5~]C��랅5�v>�����ѣ��/~Q~����{j����"����~��_�w��u��aGʇ��{GS%O�j{fl-�=9y�Q��h���Y�a�����c+Aɯ�!��^�((�S}�V��������c+C7[hϞ=�W_}�7'N���cǎ�Soo�o��x�m�"��g�y�$���x㍗/]�tvjj��d2�`�KIG%�}�h�K]������SO�+��BǏ�	�I���O~�x@&.�A�p�B9�>��e����D���$Җ3�N�G�Q�<�]�̇�v���V�)U9~CrmW�j��K�i�>���v�n�_3����/�����c&��p4YT�����������'���G��K���b��xvt�ѕn�������Ŋ�r��I��� ��Sz��p��;� ����\�ˇ��;����o��o�}Ms��ٹ�a,h���z�A�4�����Pɧ-��4ݚ�ێi�ry��j����(0�`gCm�6�����_��ւ��o����n��ܣ�>�w<�C���wFx�y�ߏ,--9�A���eS��z�O�	�R�6 5H�<x��?��g��{ｷ�PzJ�≛�%E*�P�QT�R-6�Q��Fk�E���*-���PI3j��z�JA�����:�J���I:�l�8W"��z��x'�+٪ޏ�ԿUb?S;pڎ�w7J�E�N{�=�wnmt����흫힯�m>�����v܍�V�/΍��Y,����@��������>Ў���_����>����zF�
��z}���z6��{=�5?W�|,+1Yp��^��/��p~��Z�JI	�>}��[�?�����?g�2
^p��-�]X7@Bt-jd�4�^�\�"�M ���_�'�x��R���Q�sa�`hU�]{�և��[g܊�'5(�Ժ����m��{}A_z����
X��F�g��2>���P%!v&��|V���)��,y�Y��ŷ���G�T��ǺC|ծS�$�؝y饗�����sSSSÝ��%&�@�nך~��� t�� ���i��W���eFe�X��.^-�;v?WoC+������2���'�ͅ��T�'yVk���+�ia��Z�$d�3� :���*��S��2e%T�4��];���Z���v�ۧ�������k �Z�obb�����~����R��&�z5�k=�K��ꖅJ0��@V��{�,��T]6�&_ȗ����n�;j@*ah��Ѯ5�T���L�4�>6�Jg\M. ׺�f%X^�B{�$D��Qk�J���0�H&�Vpw+�_��� c>Z���B��n�r�T�ɐN�gϞ}�����n߾�=::Z�D"�z7[Rņ���ִx�rK.�Pp� x;����Kw=*^��q �R͜^�N�Z��x;��{���U�Y�ٚ�fο��Z�f?�Z��g�@o[U)c-�3vj��}�JF����L�5��z$P�gl�q��W*��=^����F��Fk���FǓ�x�]�J1�5��d�۞�����Z+��F����6_�B3 ky���L#����چ]���Y���ߵP-FĽ698B#t�{�	�r9�=M522�qoo��+W��c�����ێ+��x�Mo�brъɸ��������E=@��6bw��!��n$>|���j��q��2���j4��7!+�ov+��q[���ulUu���RA�C*����{��Bݾ����Yh*��>H=ЋT�b?0�h�!aS��FX,�*��H5e>����`{y��Ш���VK��;�i��|�Z-Y�����'>����B$���	��B<�7+\���l8�$��7�4�	Q�C/2,eCpf㮛�z�`����>|ذ�t�%B�F�irw�ZQ�=6{~����"�n�p��mWc�>�����q��d'l��PQs��J|���#�D�K%W�����:-Ië�Y��^�*���jM:�VNɇ]Q�Y�x�������'ܭ&��i�վ���E9�[��V3�ڍfc$j�����u�Zy��h7A�����x���i������]�c�=�v���m�����g{C�ޖ��U�w>�e�{mh�A�IoJ�)��*�-�Q�X@b��O?�tL���I,�%J��ޮ/^	M[4zBM�w��-Z\\���J�oJ�V�>|���Ç>Z�5�X�3�0a	����ΞXZ^�;>�H8���Z"��
��b]�t�.\�@�>��ȱ����O>|���Ç>|���|����������wOLOO �<ÛД�^��8�OU?�V1������������z�!�5Ύ|��Ç>|����G� =ך7��A�GC&�������  ��-L[�#���@�UB2_�)����k�� 7�O�S�����OKՂI����:3��)�4�=l�^���j��z�\{a�s�9�7��L������(P�N��-֐dRcA��6��X+i�7f����f�j4۞��`k�>P���z���h4)@�5�.h���!͠��z��Z��T�*4.u��m���T�]1p�F�u�j�4:�z�����-kQ)&u��o�\.�x�:����ѹdnnn�/��/���[o��c��x��m�u����bU���T�����hvv�^{�5�����HC��WN�����h�=��NE���
4��a'���ҊD��V ޭ���� �M��4�*7Zxr��6�6#�[	�,L��&0�� �B����{����?�}�H?��%s�����< ��N�wtt���o�M���w����i�޽E�����'!kc����r���^��������cb���J7>��X<����?l��mH���k�Y/}���pk�I�*�����CWz�����?�������C=��דz�FK�z�)t�^���O~"A���J�N����+|�N����FЛj��?o�	o�>�hv�m��&x= �޷��=Dv��N�|��%^<��wH�K�bYŤa�D�țo����^{��Ν{���+�z���͒�i���A<p����433C(�I��?�y��?��3�Gn��+�����c�S���[bѬZ��y����>�u�n�.@��*�h`"V�l�t ��	iaW�\pc���pp��c�p������<摣�L�wv%�`7ys�=_ ��o��Y��=��4�:����6x]�L̿6*i���:;���7w�ߣaV9�{���F�=5��SU-F�Q�v���6�<�Z ��|��C�b=��������;^6�Ry#�u}��p�`[���^�@�^����Fǔ8��i�Z�~��iZ���Z���������!�ṱ�����vw����<�g�g_�7^�u� �[R�"\ϣ�
�X���K-�$/tc8)Ȉ.�X GFF�3 "?���׿�5�9s��?.�,���Q;�G-eg@`��v�{,���q|w�� Ƣ&1�	�#ֱ�}Mqm/���};C�=^�h��?�g�X�|��a>o��j	1v��ݾ��Mo����'��f�w��E��?(�Y�|� ��P�\ �q�->�S�:����m"b�(���5���hŮ�fBǁ�(�+����߭���c�Q��hr�H$RZ^^vx��---=4==}�����\�իW�;�������?�䓇:::����w�q���N�����%D���8^�Լ�`Nx�o��z�-I�	
n췿�-MMMQWWת]{��l4Z�w�h&Ӌ�)񱹀����x'�0�!���qVϠ������u�rb$��X���8��z���/ms���?�Vo�» T��{g��{��u/�� ���i������]��?��^#de���Wt�PC ^�JDD�_t}��%k��D= ��BQ��=����a��Oc�Ë	��˗|������2f���^&"�?������;�W*��T�^�FKM�h�|J��^a��X��1���/�Ӈ~����{��N��h�-[=M���O��Û*4Pr�,�
A�����L&U�����3I�������c�b����sXX�k��ݘ,Qw��i�.��əa_gQ���)@:D�]m�FfR4xW�)*d�����0�E�/�
��l@�)�V]�V��J+�z��56t�F�Z*���,�O�r�����t�ß���6�As���\����*�R�Q$D�"`�_����"�u�
�'�W�hGT�z�I)��ק'��/�ל�c�{���i�M"˂�)�N�k9}����Qӣǩ1����w����˗� }D�%/�����1�JK{��<g�x�`�F;�8��+#莗���[���u��opU�q/�d�m��̛�����2�Fy~��U=m%sn��vWq��Y�c��m����o߾�я~�@<?��ӓ�������Hl����p"@�䅒�M��N��sqs��տ�����w��8P-;Ȉ�^��8�e��z�чh�{�]�ˡ�R|���P����J0��vjf�-X2Kg�� �R�q����2�,�'�h9�,]z%)��B�Q��j�ٕ]�u]H�.۱X'�����ɋѮ	޴�M.��B[����e������R�_7:�\&Ka��Pķ S6���0����-,P���Tf�V�i6L�y�R�(�]�I0%�c��p{vw�Pow�t����6���]�l��ED
�9�E�F��5�-�ל/�����c��-3f�.�%�(�H�g���5��u �iz�6���1�;y��Ǻ�����
H*��$Lv�!~��.��><�a���A��c����I��e�p������'���B�g� ;�G�?�PԤ�����c����t:i+�)�ٍ�&��f���,�H|�ߦ#�-<��Θ�8�x��v;�h����W���~���θ��ZEB���y���4ma��gG,"������w�ͼ��F��i���R���`>9�����ޱq�g
�����kt�8��3�JAn/�[Jb�e�s�(V���.��!�9n��L.M]laL�c9�v�S*��y5Ii�C����,1'�-:���t�D֙eR�N&in�	}�@1�H����K]<�v���y��d��7�0��'s����<�J�=[mr���ϣј���m���\d��J)����l���T*�����8�?�r�r��l�z$W��R���Wo��	����^�;����m��N�Nwy�6٦��'��z��a�%���[���7�(]d#�#B�n�36B&���Aw��tL ��3L�����������t{�&`I�(�
a�.f�H���5��w�	��z�{�[�:��Q6�L�Y	�*8�N�lL�4;3Gs��b`b�����iht�F����x/����qy�c<��L�s�t��E��z�&�t��m�����a�����K�����%ڔQ��7�R�)(�RĎ-H dE�x�lLNNNʳ�nn����9q=z��`ts?�A���6�4=5C��Kt�Ktk�6�,�SOW7�۳��y�Y�����` �F��1/�Q[-�,��p���Ͽh���p4�n`�I0�π@v�5OMO���-g���$u߁�t��h||��z���Ʃ3�!��7R�	63tkr�&�_�.�����	������>���⻐�$��ܘ$Y�&���i�%�yAJ��s2��%لH%��.��6�/�� ������}G�СCL����I�bP����ͳ�=��$A��\�k׮���"�.ϲ��X7�S����s{Fy�f��t��Wm���P�����cI�{�Rh�1�x���F���4-%�:���C�>~��P����U;�.
�<�b�15}��j���m>��<]�|��������x�32ʤ$..�,.ϝ8"�>���E�Ϭ�:���ӛ�s�[A^� B�X5����Y�bju�L��7�U��5�>VC����� �
<w4�X;aDb���IJ��өc���?D�N��=�+�c�պ$@2$F)�Ew��B�-.,���1uQb�.�!q��y62{���'�{a�c��*���X���+R,��|� G�F�\����={��g�����}���OQ2�`�'�jm��e�6��&g��w?��C33�t�����	�c#3b�>�"��x�6��,���͉�:�A�3A�����I!RQ6�z�=���t��AQ=��s���ـ�dVr�N�izz�.~z��}�=��w��ǟ~@��C��X;^��6œ���z��`4x��t�|���樫��V�9�W�⩀4/�ɲax������}�;L{�`c;됝hx?�=��^7xS�Ʉ��9&.��;'�ߏ?��nLޠ��&����GE��6�{�EY�e'��؉��q���c60"L�
L�a,L޼!���=r�,=���t��Ac�1P�C�נhdGpǢ-�S�=���+������MMM�ECCC�MtB���@�y7�H�GmN�z�*0)��DN�	@@���&�U@<L���&��CO=��>��1�>���]&E׃�Rؕ���,�/�e& ׮\�����6���}����%!w�׸�f�+<Os;�s�$��#>ք��H�����-]9�fT4I���ڱy^Y��j�zj]X�x;>�Y�E9`t�؁u��]`!�L�oޤXW'�s�	��K/��#��������Tb��â��O@
 �>���`��ll>|��:� �a���wٸ��c�ͯ�e2r�FGF�S ������0�
�̰��	�>o���|j�z��O~���=��cb@`gv�����ۚ�&��e�vE*228D1&G��G<CO<���?���y�4���0�T�[dX��#��Ÿ+�a��;�0��?N�=�=��������i�����L����#W�Z`�{g����H=x� =��z�׿����_��G� _�� a�F��U�N�v���?< 
1�!�����!�㶉2� ��|�2�[�^|�%����=ǎQGgTdz�pT®3���K�����aCtp�(=�̓����������� l�F��8s�s/��S�g�����,c���LP:H���q�	�ɓǙ���^�b����\��L�����������}���<N�>���7��}H�������'�rq3�I j�c���#Ή��\>#�4�P�d�[\^�>r��/F�<�9���'�������	�T�	l>[� ��@Hfo�Ɇ�yC#c��	�/����w��%����ԵI:w�3�7q@2t�-����-񵀢�v���E�*$��L_���oM^aK����L��Y�������õ��ʳ��`������v�6�ː��e�w��9l$e��ɕ$�9�������'���={��/����7�]NQ��q~=��c��6j�I@h���l�?�����<r��v���g�����u��8p�\T��ȉ�\Y#����q��Τ���uZ���������-z���)�F���ݸ8%J!�A�B,a΂{6�2��S9ʮd)�]� R�:l�Jt��!��N���������C��/~AKKt`�����N	���hL��j������<3����$~��slX^����ګ��ll���4�d~�
�<���l�1�C�b\
|LA�!Je3ܮ���t@�K����/�@��)���F��k�􈕙��oLzE��X$�;OL��>�\�al�[d�`� �	��l�
�k��Z��c���������BT0N��,�ت-����0���EןG܊�o�wįg٨L����<~�I��=��c����������wlB$�s�N�3�\Zvc��?z?�AS��n�+LPA��������<�QC��"������tQ�/=
�a�
�I%���1�at@���_�=����w�K���7:�S�_9���~	�H$���sW�l�V�aCMee�Ը9�VsŬ�RB|i�<י�����������~��}�Y黐�a�C_��LL�}ݱ���D_������<���ӹK�|��s���}ab��z����������ʥ����/�bC����V(���o�;n4��VOZ�9x��x�}�v6�V�����lx��Y+;����<A�ǩ�=h��qx���	������3� -2/������"=��󲳛)�i�����#*�!}��?4"��*���1�.fC\��l���d$ ;�����t��q����O�~�|N%]�l���;?N��
6��f#sz~��nߤP<L�����瞒x���"����FxW/���.?�u���Q�%�7®`�xF��Ē V (6st��a����?�X���?�%6�-��p�Za�}���S�|�����(�<O{�/����+��4��䍲4�W��C"�!���R^��LX�LF²#��<�Bŕ<-�g�����{��'���������R�z��O�N&6�Lvյ�D�]lL���"o�+�v�%9��|��9d2�?�mq��I������׾�5�w��ɔ�?Q~V�}�X���DE���p�����4�.�O97�c��{ｴo�~:�F���Gtm�:�So_9Y���;� v*V���V$F�	޳s�t��-����7�A/����`	�z��K�ē�>"<S��Mc�.&�)?Qg8F]]��LJ�H�n'Ҕ��H	6G����7��_���1	����-�7�%��vB3a
�O�_x�� ��KA�`W=�����?IL�ɂ�(�cu0��c�+��SJQ�c����s<'_�|�n�L�}�O{�G%��+_{������K4>¯�-o�Z�]����6Gs��Z������u0@V	贳l:q�^����'c� �,M^�F���w����gh(>H}�>ZN,Kv"+��=�yE:c$Y����p�t ��1@?������|G�Y0��	�����Jn.���A�l^���<}v�3:x�Az���W���w�q5GW�^��n����P��f�H�::bb�#�!��FA`.v��E6��(�b]"w��~�FF������x:�����Q��8H���i%$�_�
sӳ3��W�>6���ͯ��ӧe����K�����!���h���Z��)�̑�/JPW�\�BE���
���#�)������C�N=�� }ﵿ������*����QWG'--,
�������n�4Ut�.9�����[�$��=�0G3LR��(��ʗ��_���1�f)TG��0QE(RY�؄ < �	
K��<�E�DC���㔀��h��-�n����/0����/�����	�2r�	��� ��9j}ޓV�1R/3AF� �g����_������)Q(ɳ�4�٠��W��-]`r�MQ�����C�	sS?�p!,�Ē|��G������(�<y���1I�ћ��:]�v�L��
3��@#iq��c�{���@����pW�\����K/�D_��Whρ}2���B�������4^�,3Q '���c��z:�<~�����/�k*&Sy�����c�R2������$pbt�"LD� ���������[Q���������NC���� �U��A6��z�Y:~�^ʇ�vэk�����o}���tRz	�9��@�I�Χ���EY�.}&cҋJ�;��`�Μ9#������K�:2��V���Z�F��
�+��D�`�֬YE��]�u�����_|����W%�.�}��9ZI.�^�G��(��pn%/5,`���Z�_bÇۓ��|�(�HOP���T2-ށ\�l� �q"����g�fc�@��5ъC~�����wۣ�5I?�*M�����$w�~�i��7^�Ç�n��?�xw�F��)C2�aB�A�R��G�i/-�Q �P0o���9�������#��;A�K�4u���h���o����_�N7�n	AV-����P��C�_h�7$�H?Ɛ�<����j�������o~�r�)\�YI3��+��Q&��|!�SR��s\J��P�|,��킫�G�2�[���x�{���K�Q���C�܋�G!�G�����t��!v��%)2�����PP��ڈW��WH�p��>r�����t߽H:L�x< Q���6�(^��?�}�#�$R��uؠ���VO_/�+�gl�����{��ޅ}� �౽���?��x�~�����e��	�hH�� ���@�a��L�t��5!`�|�e��׿.��Z�(�0AI���$_ȺsRTj�dSY
u�(R�D5��9�R�$�{�z�o���F?�u��>�$����M�ȓ��u�����MI����"�$���Ç�2J�^H(�9���ȽPC`U��5>[�ZT�����ݚ��/jipk=�ήNѠ/�͈ny��'F�������(UX�P��ޛ����	����O='�#�b�Iv.��/��D�P���̮4�0�U	KPvy��;d1���M�9D_��t��%��q��9F�l��g2�����SK�^)Ŭ��ꮪЛ����qq�29Q��<�=���i1��[�W.^�[&�đ�tl���h�a'+v�TD�����b�H5l6�C�����d�n/6��F6��ҫ�����}Oڨ������7�*y{4:�E�c�d���<�_`��e������N�3/>C'�����ӏ?y�x��������P4���,��A�ĄT�����T�a60AĢM]R�	 �z����ѷ����_g�ܻP�;I�l̦s�Sl�HŰr��Rs$��(�� �9ʆv�����牧��W_���ln09�ǘ��1�.����ྐU-ș�0�Q��M�����Fz)�#dw (%H;��ח������x�^bC���ҭ���C0M����Ʃ#��H_��6ގ�$&Y�'sv~N�͑��[���8~��$���ƨ��L�[���0/�O�qlB sd�����D�o ����+��tَ@��?y?�xL�����3A�<��g���I:��
�1G�;L2n{��+�lv~/ș ��/��k�۸}{F�v�}�Q��׾��c���M���r&�9�Q�����:�+�T��(�*q<�r��F�����}c���g���}����g�� ��R<LG����2}��{tc�6Ő
��^�\[�ةp�h�עh��oF��n11���[������Pk�Y�MK_��W*���{��U�/��pɍ#_WȮ��?1�� *ӜؙLZ2�,'��o��N?� �<}�:{c�E�8���i�����oӡ	&&���;l8�L�1,��ʢR�ح1b�	��3���YxBN�d���g�G?��/����^y�. �j������\Ys���s��>��Yz��p{t���'���z�&F���ǈMg1HsI��A������P��	���(Ea=�B���H,�����W����WI���PJ���bh�wRt��u����ګt��cbl���{�4=Ggx��!*��H$$0�x�6�w\	L ��S��v45Otq(W;��EF��,J��ltO��ӗ��*ݺ1Iׯ_��~i�n+3�<+H�Ҵ���������[�����"���������a�0bH��,��1��*�ҝE� I+�Ox�����x�2�yX ��cO<N����C7oߢ�Q����ē����"���9�L
�	�G��o�O��N?��x��	�Y���hnwW2���*
�-D���I�������;~��.���I/�e�D��܋����4��%>_��N�������ـ��J�$��C=D�'�3�J�@��9S0!SB�D��/�ߗ�	�D2^B�7$}����^#x�m�c�R���7�X�sO<%2����8��IP�.��D�&'i����Һ��Ԓ���^��b(kr?��Q��Bw' �H�Vx�*P�;F���c'���ȈdL���w���9Y܎�G<��88F��.��
$��2)�T�����.vJ������������ =x�Az�ͷ��ի���	����0�w�.�d�%#��k�@5�4O�c��#g��'.Z�T"I���_2�
ө��kO�Ҧrs�>��sJ&���^#��]a�28!�*����Jr8D�1�2��h�����q���)�G`tiA� ���� `7�C��򚳏=�i&�!��ϲ�m�����H$�=�b�"
��� �n�'����%��8��DDvc�Д���d�
3�`Ғ.H�_W�N;NG�����Mӳ�E�ʍ$ޡ����̨W��Bxq��hpdX2;a�\����v��b�	Hܐ�b��Ga�T�N��NB�ݺ#�x�c��������<��4<2H�:Eo�˛4Ǆh�gH$}�γ�˭Na�靿Q /��S��6���D9�\&Nq�ܱd7Y�&���Y��\1�\�n&zǏ��7���ޣSg���Mǎ�cG���/��A��<>8{k%jZ��|�|�(B�k~��^���q1�;,�l���y��$�P�$Q����I!��o:�_�ylW0s���#���9��1E�/_���LJ���K�L�fnNӵ�╂7R���B:䁲\,�+���۠64<�O���" Ɨ��<!>��`4i�����\�l>���x_\��.J-%�_��b�(=��#��oqi��.)W��}S}T�x3��CttS���(�Rpݟ�������O/]����}hJ��8n�*z�����@��
�:u��#A	(=�
ݺ9E��FFd������r{��c�c�ˍ�i
����Z	�X�#���nSW������E��;G��96vG�C�n �0R��d�4�4G'8I�<��I'�)&�W����K+��A>T4�����[,�n�K_!��mP	Ќ�A�ņZ��#�A���e��Ԓ�6u�����`O�1�a�I	�֓3S�<(�;��Q=�����2t��`3��7;� ���K������:�M��4�,ȷ�m���sG�Ğ�1���y���s�Ӟ=�t��������y��1n�[ago] I\�@@� "d�>!��_|Q~_�qU�9��P��!C��k_�Z0�@�BR���C^��$F)N���)2�}z�:v���;����:s���N���%~6�$V˘����y���p��#���O�/�w�F?���r��;�rY�a
䥮P���	HA>�IZ�����0Y$y��'���?�+�/��#�$���I�����E����_��� �y���v���P��^�5	/�A^0n���^[�e���K��׺�e竡ݚ�Fc�=�޳V���As����>>��@O䷓�%*@�����BG�K��y��,g�����?�G镬	�����.?�j��nuH4�h
J
J,�ؽ���!��Mˮw�?g2 A��k<}��#_���,3c�J&����t���~;B�P�Ć0	���MY���Gh����	II��蓏����0��>*H���=zW�e �8#�8��K$Y�`T�W@V%>?v�3���@��I6��I���O>��DB��H�
^���1���B:�����y�[A�����y���O>�����_�d�B}����$�	8�#��ib�3��=)�M�$�C^Cl�6#�X?��||��3�ƛo҇�}_�����*�o�T�9j�V�c$���e&_��l���'����Ϙ0C�Gv"T��d�]�]�,uA�9 �&����.��� =�H],��O�������݆z����KllwJ�CGPwwݞ��XFx�����mr�����Q������m����/���O��¬�� �B+��7��G��`�p:���ڼ�)B̘�^��5C���a,��"�
G�9B�&��y&!��
������|���.��J��`ɜF�5D�30ixx��ϝ�D���R�2�Ġ�E|I�=�a2f9����C�'�������N�� ug�}
�e��e�d`J�	��~?S�с:~�0ݸ>I��%fr�j鈓���%V'�K
i���\%Ee~��Ɖ�ض�c'����fŘ��rֺ/*�	i%Tm�sj���zU�9��V��z= 5�8>�������0�{���g�_�XWu�tIP�͛7EV�bgH�Z�iPx;@�8~'3�򤀝{�˸e2RZm�o� >/��c�Eb/�T�v�<�\��F
����vK�"0��e^�M���;0!��cw�:���W�ѱ�(�6��H����-��*��'01݊ڐ����v*��.�f������:� o��]�t����hhp�Z��I9L�q&����Y���'䒭�W��l���A��*	���]�`I�/�����\�y��K��;�b�=7��ȇ\�<�P��.-��۷h���t/��>�H�]�x�nB�l���w��Y�L��ߐAR�Zȼ4�8O3�3F%f�a�Ig�����~ȧ�	�J&���G_2������!�� ��ڎ?�suw�H�ù�۴b�:��y��?bҗ�6���f7l@�Q �XR��"��n%�"���=�LȞc��Q�[v�4�w�:�~�=(���] �E��u1T��C�r��-�QIH'Xތ#�n
�
�\,�-R��5d{B����ct��R4��#FQ�Wy&��iZmEGA�᡹�ޓRdDC
p������E#���`�V65�A���#� �r��B.+�A[��y�x�P�ՉDE�Y��=����˗.�ѓǨ��C<�H����+Ɍ�m�cB�]��iׂ܃�`�{A��XKb@�|�إH$�e�G͂xo\v�0���H��4ϋ9��LN�����&�9 ;���uL,�p� �PY��1�����HUޢ1�p�T2E���t��Y��o~'Y��rCrM�Lk�i[���� m�s��SW<.�cqjjJ����\I�5�0r�gxG�R��X��V�J�R��T*��ø��d�*�g1�(�	a�\�zE�A��<�Z*a/$ RtP2x94�gDvP#���>;3C]����2Ғb�-9�~`j^�7�RA<:(���"@Z`ȯ" B��(��7�Ǐ�s�Gi.�(��w�z���i��M1h�i�����z7b	y,t��}��!�y���N���������3��J���=♅��x��4���,`����L�Ȼ�� O@��^O�[�!¸��l�'ﻗ.��Ƥh��z�l�F��8���R���>Y\�=G�8b���߀��B�J��T��Z8�Xi���Ȕ̿#w�����zf\`��� �=�7@7�oR2�B]��4�؜޾n�NN˳C�����-��3vd�ߨ����c'NH�h�& ���	tU	x�Q��z��8��hDR���:"L�;\Y�.��b��BI���[6-�2���@���7����,`|Nd���Jj1ń$)m�6A�eW2e�H;ƒ���ݮB�E@����"��*�l�����+���V���ŀ.8RhZ*����e>+;��4��X���]��8�Ɔ��)��1(@^����8q����;��=<<,ޏ�H��@w�a�γ� ���8���H�P쬧�)	G�xW\Hh�i7Mj8L�
㡘�  k!IDAT�TA�ʱn�����Ff�H�`��qcE�b�d;~�	���R�C���WA�h�N�[���=�i�Qgw'�dC�xjGa�*u�P$#�n�¨�z%!�W��Wd��)J5�OH���U�f�mRފ�����cBa>�_������Q:r��ܸ-��΁�[٥��j=��E7!��7J���P2�}��z��
6����Z�!�3Y�B��{+	A 1 {�H��X�JE����7�W�i�n&�C47?K�T���i���4����'���]4l����؉T*`�l��]YIK���&��.��ⴐ!�dS�[o�{a�����	f�+$�?̜�����2�ŋ�8#o�5��)�'�RHݸ/���˓W @࿥�����������	�,g$n�w�#ٖ�w��s�&���4's��G$~G6u	����ِ��	�O�q��$m��$a��H�W����>ᘍ�����}����A��rl�@�
92��=1�B���ă8�]mX�hv��7���X���d�9|�;l��ll��͕��OY�n�{���vw�v�|T:�]��hu��� )�%�qsR,/�0��l p�{��r%�d)�\f#'F�p���~��D�T�Fv���g���+�)���[��w($��0$�E(�� ����@.�/ʹeg��F��8���}z��UK2v:�$��]���aaЈ��.^��	f���A�}02� ��ƀ���)��L�C�3�r�Yإ ]GL�rJ���#ƤS4}iVQ��L<���eK+t��=4z`����r��;����p�O�6���/���h	6.���;8!��J�n/L��5j9 6ce!	�E`��Q	c�	�� 3aW~������9#Y��V������d$�Kԉ��B�x� �Ӎ�[B��?@gN���~������� U%!;�`T���d���j�9�jt���G��8�IС��򳘠6���g��tƻ�x,��,�$�p=m���!	���9P��,�wz|��]2� ��(<=H���\jA�g��ؔ�x��s�p�Sk�#Z��O_��$�v�܉9t��)�{!�E"�H���|�(�eG�1��r�����/$�d����!�<`JjǄ��p�9�{�6 �R/Ddk1�1��u�J͙l6I]��m�2)�S+��z>�hdl�.}r�2���]CҞ��YW5޲^��i��&��_OdV(�Iѡ����7@�÷oMJ�z����IN��8�?Q����� Ys""�E�B���@9�W@fP����B
q&��/�����\JR���͖�Ɉ�ar�c2�>��y�VUH_��;;��l�6�ިd�y_�B���]�ڙ%�h���4��i�.�jG>�&0�>~ી���-\��~c(��Y�Hz^H�	.��zn]���؀�`$W�"q��f�2F��0
w���H��	�}�K���&��4;�-L��Y�dK�1�j�c#m����K�4~����6�TE$��)g#3�@Pd���!Mb��$�F�7�#%$����6�~d7��Ca����<��:�������D�u	H� )���$)W�-C�54�;��G��ۏ�yDѨ��x�^v���|�G�n4�B�_�S��hb��&F4���K'��h�������J�\�-�g�F�CYVW4��n��5�A�1�3
��"w����T�(����ޮ�K*�30 ;�Z�1�����}��fQ3�߱�)D����,�1�o^S>W������l2]ydÄ�K��Nvl�T�N �類&̾��V�����$I�IVP��^1��c�*d=�.��e�?c�#d>/"(l�J�``�t�� wx�J�G�g \XJ�5�i�fS{K��ҝ.E7�s�5$l@f=l��&R�L����X�������UH_'�u�%�r=!W;f�v%�N�σ�ƹr�`Ҟ�<�ISF�rNj�˜"#+�^W����>�n�N&!��C�6WB�iД���gb6�b؛���;���S���>�*���:t�#�0�4@�Fr�^�u>��#��g#�v����Ē���hv�Py�+�K��Y2u$E1��%#_^<6AJd�(��D�l�]|6T)MPt����E���ͮ��b�`�}�)���00�S�$Nj��
�Y(]HK��������'�����O�O�B5�����Ԫ�T��DQH�<(R����`����B�
A"�v����v�dV��'�i�	+���RD��2*�i��n���H�� NghpHw!q!#�+I]�� �n�u�MW�sSYr�D�XO��f�i~f��f(�H,���P�L@Ч@F�~�!6���yM&�Ҧ�Yxe7��J�LA>���p�����)I�g�(g3&�	/�Q!w�T�j<H,�#h�~��Q�~�M�(1E�t��AЕk�Ƅ�~�x/l>����%�����IBk�<��|�LԃE&/)�]�7Y��y��?�����M�TB�Hv�Hd��+ �,Ǥ�ƿ��uǻ)���ȭH,�Ox6$K\��{�!W�����l��Qa�w�܀X��B>+sG6�G��xr�.���6���P�"�3ϻ;����w3�a2�Dɇ�����(v*	�ͣl���p�&,^X�nд����YJ,���u�ٸ�J�<�]LxI
����cQ�b��_cH(`h߾}[Λ/�dR��8]����=�w��fa��|�=��W��g���iT�$�#ȄR��[���`!!�d�6�4�qN��`pIPA:���Ȁ� Esn�N�q�$��c)�H+L@F&ƌ*�)А��0N@���µ�7R#�2�sbx�Sl$�:(��JL�45fDBc�@���17�vHH��...���oR��5�
B ��徖�M�2���i�죞�>I%dC���01&&��9C��LM%<�N�EB�-�� ,�3��i66@+���J.1W��nH�`t���6��M$Ҧ  �z�q���8����O%^�泋R 2��!)��"�Yq�D�ȷ�M�v@v�!I��|c$����H1RN�*�I7~D�֪g	}ƺud�x�3�����4!Ƨl`��i�@��ya>aRL�ҕ���t�%�M
r?�慉�)���m޼�x$m q@�̥�E���@  �TM=�̈́g��E{ �WWGEy~F����,ݘ�!}�-�o��:n��d ��M�ߒ~�3�=��t��/כ|��Ç�F�&qw��R�u�c����4�y��]��>6�㥩/]�
p���Ë*��q6h���i��r��Є��I�iR�jP:�vKb6:�x�g/	^˻�&#��#��ѐ�g��,�*ː�RB�J��ķP�Md	-r���Ƈ!�\IPo� ��3F�~�	����B�Hb�ꖅ]�S�KR�0�̬�|�6�HO�!a��9����n�e��8�0;ܶ���I���b���H95,$&b�Ȏ��oM��*!���p��`|�q�ˁ�1d��{�cTʖ(:�:1HÚ�}r�Ҕγl(� E�1�BA\sI4�}�&FH�9�`J�s���瀝�@4 z��W%.�oxH�1C<�r} ���B�#��]wG�W�}�wyH�����6(�7�3@}}�(tecZ�B�g���>��E�����Ѹ��$�m���r�k�9���LZeB8K�M�cwG��L�u���x-�]�8��܌����`�k�rI� ��&��E"��_���A�����
���y }�4��BP(��py��R�����DI��@,���D�2NF2�e���	�sȻ$p$UoP���)[U�ц�k:Fƙ�~r
K�o�W2�Ţh�����}<T��&	��(��q2op�>t����*S��&
�[����2���>���o<a.�N�*
�65�VR˲Y��W�|���&��s޿�ث]��ᵮ����F��^Ȯ�f�!�plm()�w!�F�Ͳ�Z*}5v(�!q��-����x�JA)�%��0@x�������HBV"�K2� ���8�0�$>�K&���Dr�ȍ���x�u��U@A2Ջ���Z�Ԕdnl��)�!Wʊ�+)h�<��؁���$$���-�9��:|S�n"�V�VO#9q�z�Y��0q\yZA��xY�n�
I������^\^2������WB`dA&Q8�8����/��b�$�<bR	$���GB�`P��������Q��}<N<k솇ـ�b4�4G�������R��G
���-�A��Wm2�g&�5o�LP�K��E��e����|����=�ŸvFi��ܱ���2dTbC$�S�#�=&i�}��%�X-���7�D�l��!��dV���3|L��%���?���"d�Tm���~#y_|�x A�5���qR������Ɖ�Ƚ�m ��5>�8��<�E8�+KK�
�ی�g8��l���)��do�����7�=*��b;�Hٌܩ��6j@���
��:Q����"<�J�] P&`h�$�*3s�&f}n�ظ��Ř���AA��\A����
y�,rۣ�XR �����)f�H2���	o�W=�`#sC-������x�L���h=��"FYc�`̈́fZ
��)�c�����t�W�_���!�����.B�e��WaD���,� ��%#XT;%�aEޗXn���^����l��d%�U��Kw���CN���E�Bp0��4�G'cŽNف���KYc�@k���l����62����������I��>H�6��K�$Y�	]YZ)�P8�H�D�ņ��e !ɛ c!al�a�;	��hzzF�nvu�İ®�T�/�zm:*Y��L����K_o?<p�>��3�r�2����2&3O��vvKKɭ콲bbA��a|$+�[���8C�!�$D��͛t��u�w�^6>gff�📤0�%wBiu�n��+k���A�!	����Ί��R�H?E���'ә�h�����^y���S�r�I��E���b�y#��������d��d��H1�=kDN$���_�D�9�w���m�Lg��Y�2wR����4v�1vR<��|͈��w>y����%g�$!��G��Uri�l@��,��!��1ΤƴzO1�A\���V�k&��a�E�
f�;����w	�ʋ@v
���Y��0�#5��G-%S�H�s3L*!�4q(���M�!�vk���6��S����0x�-�+���
N�f��µ��%�x4�����r+��ؓ� b���X>v֫ȩ���ă͖����o�D	�@J�`Е
��E0i:a�/J�N6�M���[tk~���n�P� ���wJn6,G��y&6�lF�޺sc��wP���>Z,���u�`c����Iʊ\#,^�B��4Y<4%�
�VIO��'��o��8��>x�]�93EG�� c���؃�2Ȭ��=H�`�d�1ɰ�h�����h�Axrb`�D6#�y%�<�)>�rr��0ɤW��\�����ޛ6Gr^g�'k/
[a_zߛK7I�)R=�fl��{�	_�!����r���7��������%Y^�P���^���n4Ѝ}/j_r�s2�B"Q@����>�U�%��7��<g�Rз�98�0��!	���tN�P`�'����t��ٓ'�����d����,��&�VX�<��@(\T`M�� ��Xϒ)!%�3����~�����;�����
�_X��J���|�k�R�nް�{�NK���	kCqS�/5�б!���8�����E�_�Z*��4���%X�Pe>��@�JTPd������+X@�V�X� c��4=;-3%�ڄv��s�i)�<��*k\i��="T��*����~�������K���t���e!�4�<O�HZ�^+�-����R������Z�	n^EX�d�(�B �Eby�n�ܐ�p��XK%�(���l"c�[�4.ew���v�VQUC� �Pd��7Y�bf�r���)�Qjn�PK�T�~�"(y��� Vg+������&3��b���a��,c�	�EP���*�,�����^Zm��$`7s\��5,T<ж;���7��^�;��hgJ٭ ��߻s��˭թ�� �>����e�_�c��Z�����M�ok�dؼ\Aq��
�wzu���*����.��{��F�Ghln�Ν>�>����k�@͑V,���w����ڪlx�f�N��xsCW��QJ*�K����H9Ӳ�@�AƧP( ~�>�8����R��S��XWJv6��O����K"�S�̂��MONұ�'�ĉct��=�������g��i�2"Py���%3M���<9�&C\j�3�.��W����1R��k�6s�.��I�sϜ����yJ,,1��c���t*��f��k��4���Q��#��9菲�����%:z</D����Б>:y������P_Ő0����R�"��Ts���A���>���WZ���^_������xKQJ�ஃ{39;C�o\��gO�ɓ'i�����YZ�[_z���Y�Air\����jlX$-�ʤeW|@LK8(�cvz����Ĺ��/�=w����/���m�|��\�]�A,} V�x\4��BRy��f-��*�#CHK�(m��ZdXց�Xa:�R̮�<��p�	�����X��FF�2Y��߇�
U�[�ڤ���K��;��N����CL
&BP5,{kG��l�`B��$Yɺ{��ڵ��m�:�C�|��v��7�����`�<�Al��Aՙ��$�4��,�Z��F��i+��۽�w���$�K���(���(��&�������N��ߪ��sU+f���8�ZD�҇Lg�1KGN��u�F'�u��<��F��L����R�-D�ۍ��0U5r����t�%ɗ'n��+d���E�4�8Ow��Q���&~ \8�����&O�Y^�|΀(3T�4u���Fc����N�A���樓��*�g7�V�e���Sh���΂uЎ��ʔ�v�R�X��D�/���5�k�XW�uw���<}q�]>�,5A)��J��l���^��f+]d�񢝭Er�[.RY=d�M(��41�H�bT�F��߿/�}���1���'��å�q)oP>�BQ"G���t��Z]Y���Nz�����~BWn^���(u�w�F��X�]BIBKV�����x$-��EQ*��A1�L��W���3��8��S)��{�w�����U�(U�|/\J�N#��S%Ѯϲ����N�(�^�Oё��t��]8{���]���CR�Z2�ق<�>q���&`�!-�B��P�[��*�h���@I\�L�n޺AM�0�9{�"ܮ&��E�`AO�Wd�B07jv��%�j5H�������c׽(ٿ�)Z�3��f��(��J��V�����_��������cz��_��2�PRP��fa�����nA>�R�F�J[�S���tbB�cr���)�v�]|��=s��Ǆ#�J����yg��(�A c.��4i��sS�`tL��w�:��ŋ<G��{��OG����w��JP�?L�`D��e�R�CJvzw��[[)k�%�U˱���g��7\�@\;�����߹)�㧎S(���Y2�%�7Iʲ�]*X��g%i�=u�{(9rm�:�Y��ď��ivf��1I=r����Sk���?g׸1˅�V�))1� ��bi )J)��Ų��1�b�_^�q��BC����n�A�_�@3��b�͚V�g�J4�tM�y��ш�˵�y��>؉�S9��4;���*�&�U��=�*R2�Fm�6��O>bA��(�8"�	6��s4s�n��Ps(LϞ8OIlj�c�-M;o�k�	�B���I�:W��' !�j�%l%�Q2�W�{����#z��%::t���&�-�D��픨���߸�f)V�L��
�tF�����(����/��'N��ɉY����kL�^~�j�D)OQ4�6&2�;[�ce)� kO釭M�Pb�j`I�i7C����O����K�Y�|��Z��?�%zAl�ͭR�Y����EQ�a�	R�>x8F-�-TL�t��Y�����/��}�˯��#'ĕ
�%� 
%�,��u@�J`�s�ɩa�!K�d�"����W��k��k_��?{����)�X����D�B�E��C�~�ȝ�Cuq&1=�[���D��k)�l޽5b�駁Ӄ���F�}�Ez81I��˟Q,�E�/���5��u�ڣ-B�@bp� ��vmڜ]bgX8D�+���	��([�21�Y\��k�>���g�{N
�MLL���2���XȘ���U�!���f/��p�C��X�����ޗv��H"�Lo��u����z�ݟ���P�ٟ�Vy�JqMv=(?��:_3�ayXLƩ�R�ϲ�^�P6S�sk�S�t��ZL,өg���LVyl��&{nzZ��WW3bQ��l�[�K4(I!I{���J���F��{��W_���A:~t���H7��t��9�&�E����qP>X��VV+,�ޠU[Ȋ�*�5�dZ�R2?P�gŅ�>|@�L�L�N�;-Y�����;�w���ߛ��y�& p�CC�È}�u�\(���@�`��S
��)���9>�T�M�`c� ������w�Pgg��a�����~j
��ڧ����-��<I�=�Z��h���姜��5A��b��q h�$��G҄��F��?|��8u��{���ԣ	z4���f�p[0H�t�j_H���`)��K��d3Y*����̣Y�{�=�����^~�>��S0@��/��
�wvP6���0�� ha��]+̼�?�_�ˉ�N&\�XĤT"C���7�����^����9(��Q&C)&6m-��JR�~v���s1���45��R�"�J��?E��ޡ��������@�>�J_�T����1	��*��Ŭ$�Z�<HM��YŦ�'n%$d��RV���F��'�ҕ���3�����V�bxW�V��
1�Hf1s,m�h=6����<2���͹�yc��}����F�5�d�G<g^��7��-���{Wj�\z�2uDc��9&֭@���h�ߒu�_�`��0���u�J<U1���fÃ�����[â�~��%&	i�Qcb��Mz5A)���1^�="��=���͑fI�0�p�n|q����A�L��:F_z�e�ٿ��~��?����?��+Y�;>�"#X+@�疗��(�K��4_��Ob�L��x���;��(��^z��W��XR��C���d�@�Z��#�j��;� ��8�����^���#����:~�N�9-����̒I���x��Z�Rl�U��Z�A(Z�qOPB���`�����4�J3t��u�r�:��E�{��Z�//-IA�)S��b��6���ܒ5oh�R�	���a�>)ڭ���%�'˓+��+�s;4z��T��
b��s���|N�[�Vk�F5<��+�s�d]A�����#��� }��gƦi���x��ۣ���-��3c���]�q��E���<�|"L�n��� ��N�v�(qQw���1���'��ׯ1�8C,�qB�4=Cׯ\���e���%hvʹ�����C"�3��|�L�ge3��ܖaj�ё��ܾ&j�l�g_�H_|�]�"������@� E�ɋ_6�
�X��ô�� �6 &��cȢ�`>����i���������t��Q��%��gW�ƵL����e��Y�0��p]7,w�J����.<�^�݃|���)g���&�T�v���Ԙx��E�{��_�ܯ���7�F�����p���4O~У1+fHjр�LKD�)+�x�hH�O�����5���� {��z�-
G�D�����w���}2)���%F��dNEԘ�i��)��S򃁰'�����7)���Y*�E��� ���oя����_��x����e�o�5'��� ��A���y��j�C�$"(�D���;c#t�&ωT����k����(���^eY�_������t�H���U������r���ÖH+-�/�O�o4��K��9�Di��\<-)�?��G���_���oRo���ᨌ��s�x�I�/^K���w¤-�P8�9��^���i�w�n�ߥ�SG���s���fĲ�hl���)�ϰ��<�a��"�l����N���8����s���Ss0B���0?��{�=�/}���ON?��O�AgN�ŃhK��g�2�Kڌq����/�6beIf��V�I�������`bLj�`m��K֜$��[W�iqz���(�y	��inn����[a7�e�e3�v��q��(��W�^%$塚^���Ķ�7�lSSS�;-��Ʋ�hh<%����"!�Q� ljf�2!)R!L�,�V��|Nm=1j�������~����]����	:{�<�>q�7�6ZaA�p��&lz
�z!V�j���2��������o�����x�^��7(�JؼA��?��򙴶��G�v�������2GXpF��J��� y&ݼv�Bm!�y�h-�J��=��7�D7�ޤ�7h~y��b}t���l��cD$����I�Bc�n�@��Ԝ~~�᣻t��m�y��ӷ��w��c2���ss��G�R&�a�徐m��G��2�0%�Vhu>�x���,�#D�/]���+�~F�|�+���g�2	��I�ƜL��|��I&#�װ��Jt"����H���'����^�L�Ν�hG��.���O����xD�%���V�c��=$�$��=�Ԫ�2�hN�7�L��C<>�j�j���}�~��{���~Kc����s����b�B6������J;�����b��E�1�.d��~q�s���x�����бA�{493�vJ��(�5+}�!��{X�d���h�9�5`��(����R{o;zB<g"��+/I�~�￤YK�8O�]�y��h0�Ks�"�A�����%
0�_L�S*���wn���C���h��1z��������8��E!_���b4��KZs� -BV���|��Y+m�X(Pi|�g��'~D/�rY��7�������?��?�i& ���:��:�-�J����e�L�����x�[C������>�1&�����ԅ�Rf-�3x���#�{{���#._��Jg�/@}v����������\O���Ŗ�K*}[�F3,�,1���ۅ�t�Z��F�/� ��xC�Po�	b��96�f��/�R(�ޞ^�(]W5��556Is�q���'46����Q4�L��m�X�ix�3%_=jf,�Whz����)z���H���_�A��OHJN��������Y�uSKK�����䚶K���[�K��e�S�0͍�S�F���O���pvy�b--t��Y�����abn�I�,<N�LF"�6&uQI��<�K�+"P��"�Hs�.���$��+���Nѥ_��#CL�2ܿs,<ehtt�<x���ڰ�q;�{�2!����Ij.����G�89#����o����馁������L�p4=IG������� 2�����	�r���S45;CK��R��.��˗��`h�g�g%&��6�-��SW[�h��إ���Au���8�"�������Y`!wuv�����ڻP4����)Zc��F��o�A_|�9�>���E��Fx�H �,R�D'mΕ���YYb�4�&���En��I��E&��x�r,HO���;��4B�H{�Z�-�������Ք�&��`I���u����{t��/h�T?{��P������FW�?�_�G����'����z:�)��[nYH��@�UÕd�f�yݘ��d�Mt���cG�2�N����f2v��Za�������CV1�Q
ȢQO��q��q�q_�uwk'��,������;��7���b�m��~���r��n�����I�?�<��qK��A%I��&���q?'��p�<|�kԼ�����>)ЙH�J���'Ʀ�Z�x��#�d��x�@�jni��G)X�"]�Pc/pX<S
2<e�fޓ�mmm�^����Զ$
����ݽ{�<
#�\�44�4l�ג�j���7S��n"�+L����F���*�mko#���I�|��B�K� ;33-��",d�����f�fm�,@ �����k�>tb�^x�Ej�l�\�$�����}���`ᴻ�K�1X>|v������EMi?$03�t*G��e2�D�f?=�5JG�wh��a/MLM�`o;y�z��hfr��e���
��P���Z�[%��Z��n�G�7�l>��z����ԙ�b=�{��l����k7)�m<rĪ�R�K��j��5Ĭ���H����IZ��K��C�a5C͋��5E��D��׿B�Sst�o�3v_��|��`+,����w�� �b!G]C��ܥg��+��Hż����*�;;5CS���Z\�$:���[Y��⦷1ճ�H����6��4=>C=SB�$A@G��Gۢ��7�L��y�[7�i|�!�����:��]�� �@�?�� h��Gy޽��+�h	��C���)Y�&�ɗ������l��~���ô�^KV��zA�1JV�nԖ �hmn�ޮnZ^��'~Jޮ�!྅�#�N'N��wJ���?������ r�h���
�#�
uu�W�W�Y�^��n�&b��Ab�V��3����h��EWKe���q����0���B�a�!�C(��536֟1d�@�G-�#L�����/���~钌��X����t��Q�q�&��A�o��1��=&	�MA+C`�$�gX?�5*�
�p�=~�(�]���Z��#�JQ���R4�,ٯ����)�/ �hba��#ɇ�4�b����5��{x�cy�b�������������7�٬��$���'*	3�
8�r��A���\�nn]}Q�0[QR�"�e�<��dqA ���So[M����'7��(�/\����)���gZ�.*C�b�(�����]���Y�Ж־�g�߇���3X�N����.����sz�'� _��3�OK�<����mA]�.��wb�1r9Kc���3D+	p�W���J���)�����\8+��@W���Qs(BG�?�O�hee�VXP^�Y�x|E�iļ�R��Z�.�����M~���+���KKqZ�����)��ﾠ�����0͂��3��ӮA���r���c�|,9~P�?CeQ�����GŹ9���e��"|�[�^�4_���#f�he5�D��N�>FCGhm-E�S�����Bj��&�X��~��Й�NK�޾^�2Y�5-�ٮ�|���9����4�ܺ�c� ��`!CjU�6�ŦT���,X�Л�[�W�Γ�2��s ��>��햠���e�{�wY����;�O�L�R�,5� (��:����c���1dI�;���)�aА���t6QwK�:;��3&�liiA��HK�YZ��{4?:K�"��)��\�cs3�IT�5�A����z�5���C� �������~!η�ޢbР���
ǘ����ma��i:A��1�S43ҾHS�YJ/�ք�ʑ�0�Z�$N���>\a�\Z�w8�������V�V)n��cjf^�?�/"�&豾V����-D�$3�®�z�v�y�N�3F����������(��<6@���Fǎ�uc�WxXY��i&�;�i�1�z������B�J�E�h��-�(�� ��'����Y�i��͐��v��h--�Ln���R�PҲ��c��[�F����#���X�}��|.�3�H$�v�ܹa& �[@x�.��?�sL@��Քi�r��LHL�U3vKB4�Z�(�4b��X#<,�����^��/nSb>Ngϝ��gOS��-\o�6�%�*����d]�!U���#���Y8ifa ��xou-N)"!�������ѯ?� ɾ�A���[cm/�j5����X+2�|[4�(8re����ĳ'Y��|S��ͤh��,,�����"hp!+�Ds������N��;��Ņ��_^Z�������������y	h���V>64��,�,;��g����(+Q0�����8�.$� !��ݻv[|�/}���R�R����y D�b�9/���(�
 D��#��'�
�iiqA����L:���C�/�)�$$$���W��A��Uס �C����J�[�E��@�̉� ���Q������$5���<�<�;�����b`�F�Z��	g�P��(�
ҋ��9��L#a6��	�tnvVNg�r|tL2)%d.�X�N��	�������	}r̛zg�*I����{ܪ&���ȸ��N?����HU�B���p�����
�U��܄u�'�G��a-��e�AP�.F�n�P|n�:��T��cbnVbA`�ho�I���띅��6v ���?b����������K_y��<s��b^��@z��)�),`��l�`��c%��e�����#�U>W��~ą,��eitdL����$	1P��� �p�J"�&�=&vZGC�I��"� ������C\�9�X��i�r���+׮]�c6#,Ş��ڡI��F�l(xe��T���kL4������-����s3 ~���ȩd���F5��%ܠ`X0@-�&�A�!٥X��%�d�-�^���<%�pX�[7n�M& +,`����.�đ	Gef)�ۋ *����|nh�A��锸���<���)�_Y�n��t��Vjjn�L<I�dV|��[#��X�}ؖR(�����V�M[�]�G�p���gD��hi��� w�h{�M2�������%)��Er/I�j��B@����ӏ>���n:v�(��V�l-0�[�Ǻ[(��[�n{^��J�t�֘\�/eE���=��Y��O����Z�f'g�� &�ko�v��Ҷ��Q��+�e�लIn�ߓ<=~�n�ܤ��I:~�Yl�F(�[�H��H�-����u
�dZu;W�+X�)Wג4?3K��o�U�!3@��5I��>�7@��]V�8`!�B�) �k�øF�=����;����v#�����47I�oO�/���d���Z���jXGQ��].�� �Y�ר���4�=,c�_�cR�����8��	!�p���dE���;Z�ʲ��G�l!��� �zH�{o�>��Z��x�nb=��I��.q�"�][O��X
Q[	
����UԊ����7�k*�9�FF��'_H�>�5s��$i5n�m��
�!����̂Z���.�k��Y���/|���}o```$�E��m	&����'���o���O?}-�L���x�^C��I���$��4wy�Z�$�O���) �4�_'q�y8E��W�����H[s9�#\��1�P����Q���w^W�qJ��
����_�M��ܧB*'�BWg
��8ݬ,?��o�Z�,��Ұ�@@�#�Qi���w���2�>w�Ξ=+E���"Q�8g��U$Z�T��`���EZ\\��YT���0���ۨa�jiN�����]��!x]bk|�_g��R��{t���Z�X{��"��!hZ�V�O�`�:'��r!x��tH���Td���|9��"LEi�-��CpF--/�������[�Rbq��=��Z�ZBQ�m�~+�0���"�K��:Zc�:9N�|ߘl�v���-�-�E��3�	����=
ǭ���%X@��2��������`tT\h`YA�:�a���D饔|��9"B?,8��F@���"�{�"#{	�K?���FB
���c�L��$-L�RܰN#sP����}V� O���MC\���)c��=73O#w����2��7U�H�C*�����l��I5r�5\6�/y��_�x&;� ���@�%�+��3�\�Z.�L�­Z^�9τ��<��2
���O���|��ϋ��7Gs�S�h��(0Pi�9%I���aB�"c�\(S�Fc|H
d��VC��.�4.--yyݸ��o�"���RXa{ٖ�`buuu��կ�{�ĉ?����O>S��P. Վ��[�[W"/�s�	�A�G�������[n�s8�b�IC>'�T�<|<1�D��y�mXX\���ajmo���	LG�@l�a;}~.ɤ%!��UH�}����&%���DkGuut��h7�JqiU�6�OV���;�	�o�����b�D)&c~�"M-�aR�M�G3����(��>A��XW��m(�A����*��[iX�H�`�f�z~jV��!����l�$O�dA$+�����K,�"���Nl�}�M���̍g<ҽ�n�1�LS"���܊�CxM�V����iin��bm�MBP�Z���p�Ij���"iB�[I
�lk�Alҫq��X�1I��֦���  �1�$�$�ԋ��i��ӦM}eT��5��58$!xpw�<�<��:��'8��[ �{��$0�/���{׷��SkU׮�S��Ww����89Fs��~E�R%S���઀,�7|F�w�&��CXWs7���&��4�vh���A��q���Q���9�V	��e�JY ��Kog�����7�mQ����k��&�+?��;~x4n�X�������<���r�r��t/�IQ%��b�]jü`�@�������{����>.�{nr��l3��27'w�N����f���F�e��Bs��䈛���VM[:��^�^��z��$W�T�l^T��ڢ��?	�4�!f�&�:s*�F�Mù԰p��ܼ�:���'���Ld��ˤu\s�Y��a?�>'k׀�mju���Kf���Z����U�R{ۏ~��R�);!��L�-��.v��*k���#s���@�.�jViV�����`d��buA��c�5�x��D���M`�=D5C/.i"�U�����綜��֔]�"�l�W��4�Ε�(�+ݾ����@�`���y�����+�-�gq| �� ����D��%3�OT��Z���J�!ר�U��������q.�oLP��^�*��6�Mg�`bcP{���^f�/�t�R�w�����I/���䯃M�_^��n�Δ�?=�կ_~����H�Xp�Ƚq��uKT���0@��-��q��O�����p�"�.�y��&ޯ\�L�L���q�ѡ�h�4������J��M-T�s�>��(�>
����Xyܖ�s���_>��"��%�Ϩa�}86}u���M���}B��������fpK�-W�q��sg��v#;��/�0�V�w�n�֚`��tJ'��d�`��1�{�L��6���舟rvs�	��Y$���K��~�/5��by7��ԥN�g���,��{5�!:�(3Tn�>(�e�����xl[�r��oе�PK �z�����/��<\����%�OʯM�+.��֙���r�b�"&5bA�^Ƴ����5���;�/S\YX���f��W�c�T����*�bu�K�D�B..���Тǉ��	�?�i[�vM��!�m���'q��Р� 
;s��G�eq4�\N-̊��}�1�\�.������*`����� ˘$�3�Li�T{:>2c\��8���)�(����3����w�Mr�c^`��OzqE������j��ٌ;l�����ĈJ!`fޥ�.e�1�Z?M�\�Y,ϒ�W�9e?�I����JQG�2�x\��CX�)J��9��!�95Z���ݐ���In��㸷�M�����݉I6����r�Q�+Q�a2+���5�;�m,���s� ҳ�l�U8��-a���KF�S��m����Β�~GG�r�6��l\<�oo��6LF���}��u���ݍ��8�/ϛ?z99���[����vۅ���.�0��>2����p���&}10�LqT�_ۣ_��n�ƔUI2�`7�G�/t�a����9I8"��VԔ�HHt���H�\\�&2xCHEzH�s?w���n>�QU���1�
�sʢ�gm��2���..?Wk�wGG�x
^�i?2j�I�a9�>S}�V���k|[Κ<�9m�9e�/\���+��R����)S�&ƃl���{�����@\���^x�U�Ht0jN��b��#��Wx�RZ0�e	��s�ߟ|ةȠ(q<c}�|��||T��	-�hN� ŭV������,��D��Dʄ�ߝ��?�+���H7:;��	��ͮ�L�"����c!�v8���(
�g����@�4^������P�Sˑ�@#���\,ޭX5
�:kiT�E)�!���j�T�C��:z���׹�9�4#��t� g�x�����[����:�q�LU�λ�����e*JT�y��u��n#B���%ʩk�F��dJDH���J���Q�Z+��~��+k���Ag�x~���[IR�WN����zp;��Wѧ��$�BR:�Z��=�̶N�̹����_գ�4~�������¼�ݬ�՞}5��O��-+$����F��|�� ���/hN{N�<B�����0ԕ\Q��i87��}�1����q0T{�b�/B3f�ڴO�Mz+�Z����o2�`9݃ٚ��l�xY�,C>
g��])�z�մ�����?R�U�u���/�F$�X%����kN*�51X!�a|�h�Ȝ[������WL�3�v��N{g�N�&���4k6R�N�ˋݥ��Jb8.9�mɵi�4�E�)c33����@�ej�gdO�A�Q�0M���?/ �ȹ�G3e�E`'�"�7dO�+Ș�߆��u�����>A������"��r��׮0�<��^V�,%U]��P�/�_�P*cu��e�k)HYw��6�>�Z��2o���w^��S=(?�e�W�G���6Z��)��b�%�/�Ғ�_��?RlK���p��̶��fb��F�}�D�&���hl�}q3��`���"z��Ӕ~Y�wQ���y�WΈ'Q���9/)o�)vV���|���%���V\;�a~(tH^^=�L���Z�?�6-xQ��y�h�[��4��z����Wq95Y�v{���S�I)B��-U�$��D��W�=rl�~�o��M��o���G?{���o�I�����:�Oz�D��d�Ll����]]�u����g�c�@*���Mx.����[�R7�
I�u�馛��7����9y��zO�b�k�f����ZJ��_y?�ljҿ��R�B��WA��lf+k�@=���ַ�h�@e%i6��6F=�3�,o��I �r�yV�귌"��l�M��]��*�c0m�U���k)r�W��,�_;|o���2��'��2`��ۭW.����9�O�СZ��4�P�O�y�:�Z<G||f�+[�']'��3d(�����:���t�x���2�c%�������)�����3/aW���֖x�5�uܡ�F8~�!9u{{;���?-��� +aa�n�ߧ��tFl�iT���9d���1G�:���q�7q�d	Ø������1]�b�P��oF1I�#��:*笝8S��g�фyp
����,��	���1�g�k��x���6���y+w%Wx*�SW����f"Tǘ:7�?=�Ps�u����y��0����q��1��+���#i//��?3y>�(��C7���ꝧ0�G]�+G��k�gJ���;0�*�7tL~"5X+i�s��"������m�y��PJ�����F��%2�3��B��	�jWD;���E��#h(�o�?}�V�#����M �����1���<n�Fi�/²������A3��v���QW�jp�K��!�,���Kr����D-璖IpPd�ݴl��g�ʦ�!�)W(�獳 %Sj-�~�4�\:9�w�LA�k����x>�����t��)y�wwXc:U��0r�c�R2c�RG��|��=!A�$y�y�w��������������1K���ݯcbK�+������;6L�M�ku�j��c���dzk?	O`��Ж�5A���)����(P��9�x�er+�Gi<�5E��r���#�X͆���\�˞��3v��<�&gK�%RM��f��T:���[l]eX:M�]�%�|�^ ��c���pv�A_�2���U�0�V+8����W-ɀ���4L��_t
�mv��t�#.�a���UK}*�溱_l����U��~k	��0>w�j�!���ޚj��.Y�h�$�y�g��$�%�E�i���0,�A�K���:��~��ӓ
W�w		T��xU�N�:P��Ð0*�iĶi�}'�~,������I	X�%0==TWW�y�H(���p�֓mpf���pfq�jӀ��;�ܪ��s/������b2q��%indA�����t�o������f�8���l���'�AH{��q�#�8�2��C۝�s>M��M����y��4�aaԍ�j��/�[�{$B�AC+/6��?)�����@�UMg�H��.�.���S�Q�&� 5Q��I�4�T����k����'!�������6�7߼p�g�ܟj�+��e�g�Y�/�܌��mt&~4`�D��tw�E,�{�>�*�D�9!Z�T�\�K`��Eg����>b���.�k�g�,L��-���<�=�AO5��[� =mw�js��7P���Q��,�.�A��،��'w�z_gg�^�?�[��R�yK��,�b|Z��w��jO�����.
WHwby�8�x��w�h�k�7+�u���ou���X�0o>m@���򳎶['$6�[\�� p9ڱ;~��4������4ͪ����|�#ךE��-�.
�5$\���J�ّx��K�v@�Y�O�&9���X@qr�o)\ŀ[�n�S��V��(Ґ�P�s�kJ7�GB�A%�:�4�C��tz����Ͼ&ZS-��	��`;���@��k6�}��&�Ƣ��v"�照�]��w��@{K����2���lM�l�S�����z)���ߌ�=F$o�Z���q��m�/��Q_/c{.�v�#��344��d�S�_٧w~6�H��yOa����D�����3c�F�vU���5�,�H��6��_�!ZLa��2�6$oa�zmi��K�#�K���i����N>�/�~N~��! �����6O�W�Y�7
�T�op̰��쥫L�a��T5�Ԟ��΁�`LV�E�ƅ�N�g�a�T�59N�M h��c(@�=�^�>�����3쏩;G���D@�T�sz-U`�K�Hw�9'�/]����)�Q�2nn�!�M�;�c�}m���(��ۋ%.jîo�&�*
�-������YQI�B�q񍅅���˃Ǳ�2���V��&E\޶�;\zl��W�p�զ�J' ��C�w��[Ӈ�4 m���Ԟ����}�[@��»a�E�.��Sў�Y��;<E���<^B���G��
�\��ε�`�br����x �~MIS��(ھϰU�ڷu��Y����XXr���.��cl���}�c/^U�T�5}�?rkN^5�.���Ҕ�hU�1�'���V�ӉV`���VC�����P��v��S��IM*�d�]�k��ewH5�F@Ϲ՝�K�6�G��զ̢����Ҵ�9��K�R�>Z��	��3�e��FC�piPK1I��#�P�6`'*�t���G
�� �j>n�Y���d+;��3�
������^a�]����xO}w��{��Ѳ���S׽G�Ӑu}��񡱪{�.�%��MBf�Y"5�O*��^/�:RM����"%�5�^���>��� �զ�|LH�����D��_A�	w\%���C�Fz��tlE���r�%D^@�Vu-�&!&��-�Y�x�?��eX��:�<�>}A�D$S.`P�Ϳ/�#>���Y��'���/�l=M7P,h~n�O���]"F�_m��������43�_����9����"'�"�����ۦ�0�(��jh� ���;VY9`'y�z�-#4x��������6~�8��.�p��'?i�]�%��Bef�_;��c'}Y�	i��7��{49��C��
U2��Q�%�U����VW� ŕ�>Xң�����{v�)�٣��*<��ۏ��F�z)��6�'��F�"��X��1����[���_�� �����kChS��H�]�Y�����q��� v�Ҷ�¬~u�+Y۟zD�Xv�cmd$	����/��ʜ�Y��Q<�L�����[�Y�
�@AAABR�z�5Z�k��`�T���<WT�$"  FG�Ok?Cu&?����/�c�:��dĕ0)ic߫��6��v����'�V��Bʃ@e_ӺXe��5k>�$�(��~#y���PF�G����mWs�3U���m�Β����y�:%��^1`ǲ2�k�-Ah�Q����g�4X��;��tU�9b���6I#��Ń��"X{���U��s�����8�t�ފۡ�h�Au���7m{YN��=%ՠ����+����Um�K/���{~�;��5�R�|s�QZ�pyV�y�"��ԚGB����W�a�&�sѭ�W�%s�ʂ�A��;^�`D�6 �PcT�^Xt6�w���k��������5����*�h[Fܩв�<��C�1�5x�pk�}� >��~<�ՀC�)3,W'�[�{�B(&���*ط$����#��_k�xb���">8��?�� �LO�=zJ�a�Z���B�%im;���mO��"���d��-�z\D���^2?}��񱢲���AB��RN���W�>hٴ���6���I�g�វzf�l���͆k����B�T�|%�A�ƕ�b�+S��������ofnhA�SB1�%>������<��Ĕ�C^��s��_<��-v��:B����r�xl0�`�j\s<��]R��@:��1F�yg�Oc  ��7c�%&��FB�����"0������`��ᗚ�Q� �G�}�0mޔ\��7y�H��c����m�~��(��7yi�0Q���������E��k4?�C��s�vg����j��BZϰ�P7!�5���X��
�P�_wU<>�<>�����cd|d�re"�A݃�d� }��<pX)������>�ne��,t�pRȭ=�+Mw�P���
�����i肩S�����B� �˥�s<MO��M��дR�X%J �����
E{>��񌼧���zb���g�GX�ν%'[.wzERE(8R0����������������vOH������ ?�fӏ���bt9Y��=�����w��.;b~�w��Ū�_�X��SHFY��p�٣�7�����rxI*����N�{�,�s�"sW&s7�����7"&�崺����V����>?�n����^�������
�|IzSS��c)G���WL�TL�d����Q��U���!���q ����$F��Fd�f�<��N��mw�`�i(To,����c�E�cG+s3�����wғ��d^�s�̷Q�	j�lI�:I�9�;#�_�7ѥ�.�3ȍ�c�@��s�	Mz�x���P���`�#V��-�3a>?���7}����XD}j�mm1�PX�L((���w���M�`� ۮ���u섦��wB��~��;3{5��8^U�&��xL9�j
X����1fܯ<V���j}s��D�ca�TȊ���`5_��u)x�fh�#�S�� "��d�v�v��|��um%dЍ�*]�Z	�3�S�<2����<���F2~0�F*��o������΢@�9�7�=��0\*�v�C�Ow{NI�����V���Y�-�ex����mcYt�i�{^e��pː�:E�@%S���B�b൱��(~<�f��o�0���seE�ba?'�c����pq}~[ǚ��j�6ɗ|f�m�"�x�֯�h�@�>U5ȉ"ne��Y�X�Ջ�!Rn�����T����	�*x��hڸQR�Ǹİl�zF�G/mY��ʽ�k���[�i
�}%aW8a�=-=��ps�*%�bR9�����,}���/�{JG�utGIc��NTfd��?>�֯��)�	����eH555����E�T�SP���Iid3[���rrr���="E��k-���3��bc�vL�	��{��y�I{~���AM�%Fo/�lCE��y�ZkF�Wy���U��_��6�h��BI��k�k��{���K��k�YK���fi�;��@h��銜��K���X��t���2t-&h�ž7�0�ϳ+��i�c�bC,=<<
�� ��'��D�E(I�ط�a���w6���	� FK���Z�`�>^^��?����������Uj�wn+KK�gqC[Ҳ��S�Q��r��|�5�n	8�� bn*[���m!�y��%���9�1	�`�<��k��Օ�:Ғsi�Ɯ��m����21�*�m�̸M[�����r�t�C��B�
�d���d�O<?tp�ǅB�Wq(P�[|8�� �2�1�b��(:���Pc�g�,�w��:��(�c���&�en➎	6��Ԕ�2G.�)��2���l�ONP�c�R�&'K��_��O�_ʿ٩����ee&AZ�y&���:pg'>��yYfQ��$�)B���z(z�@��e���F!�?�A@L(7�\��a��(����ڷ�"�.h~BI��+�_R�WޱK�Ѭ���dߩ�kdq��C@B_��:�l��F;z�i�_M-�j�#��0D(f����CS�!�y�(��'���F��~�uFG�.x��ef�0����I�8�u�~<���F��e--K��}��/����&L��ؽ���qu�2�MGMM�>�y��I9N�m�3uq��R�Ǆ�x��r>�7n<θK�ϱ�;uoY)!P����݁(l�����������綥���n��F�ϰ�=H�k"�oF�1�ף�C��b��W��%/YG�3�x�<�X��hAK�!+���]�Le4�U/u���o<�����"]N��2��<���W]s\�=2��q��ڏ�y���c8��H�i�I��.N�	��,]��lǸՖ�ߠ��A �(��ZQQQ�Z_�f���++U"�R��sߎi���~JP�5"(Zy�(�>�s`�̾!54���%L}-Q�{F��M�����s���L�o;�_���Y��<��@�j��h�b��=۫�qe�g�>]�}'���t�*t��CYh�"2�C�C�+F-���^��=�Yt�mJ��v6(�_� 5J�E{����w7��!���C4����p7���*ɞ�Z/�뽫������|������V
,v�X�x�?N�F��ʯ�R��"�U��W};���m�2�-�)��*YY�O F#��g����������xoɵ���8x�ʵ��{�Y,�J���ķ���޷�|��e��?
38�'~�g����p�������^.���N���ÇS|��,Kkd��~!��e���$k0���3E2b��ѯ���ƖA�"+�����*ܧ�4��W!�
?_E����P%3���k�Wfۮd+P��?��ۺ��"dh ��BPԽ��e�#�o�?zs�/��ܙɽ�
�Մ*�ȼf��K)����1��P��D�D�7��is[�V#����^�u�Hhx��:$اa���I��r@̻�x�#|��I_�1�>�їA�m��$�#]$�Io.�~�.�o��z�I>�c%���\�. ��R.�w0n�I(��e�����d9(˅��Gy�u[��5��oﶎ�
����h*)ڄ��=rn���]S�G�d(�7�j~R8��ψ!{i8��\���y!��eI0��R�E�<�;��!Qnc@ѹ��1��^�#�	}���u�?9��q"(A�PW�� Hۘ�s7L�Ү'd�5c��`�c�����yr��oJE��O���$(�y7����<��Ղd�n���{�lf���)4���m�C])ޮ7�1w|�5��#Ϝ��K�X�pQ�;+�A.56i����,l�:�'W�o���o�C���T%��T݆��j�v:8���xJ.����F�`��%C�R�werU��ſ0TJ<��f^>|Lf�b���?C_��[�2�}F�i�΃���Ha�q�g��R���g�cX�`����{�S�D����\���C
4�ͯh��?W�;e����/�هkC��wnG��v�X��r��VUWA�V-I�5�p�F��.�߬��6C���c^�Y���� p��힉�I�GH�����Ξ�AM"v��u�V��奻���>� .�E����	����k6�����ߊc���6�'w|M�4��\��	�(��]6��EEa�J����i��F�r)I�71���8+=����[lP�����d�pGfT�9*���P:��[��Vq{���E�u�%WQ8;���E�p.����(����ƒ^�������{6KIK�H�>�
wZr�z��N�ɶ�ð4;z�� 0�����ֵz�#��V�J�V��j"���!3��&cs=�n�	
{��ꥬA�
���a��)n(�`����=�	EI����=��޴�a�?�b��GD�w��q[�
m#�,��+7Y�br�WI�����?�9����2�`'�:F4�0ۏ ��9TZ�u������y��`��#���ಁE�t"���#�j���J�O ''7Tʩ�sN���b#��(i�e�Aq*\P����1��R!J�;(q>��Z�U�Ũ�a���q�����[����m�_��a��䟻=���%Q��Te'�	�Ÿ���%��p�x��J��w�'�U�Rl����?PK   ��X�,͓�u  sx  /   images/a2b075d1-9af0-4984-bc8d-fa1df8fcc417.jpg��uT���9��@���w�%�Cpww'@pw	������=��|g���޻�o��WU���tu���m�m�^VRF 0�wޖ_ ���i��_CBEBBDDBGAAF�D���@�����}��������=�<|||�w�DxD�x�x�y¿{�А���0�������
Gg� G�ǁC��{�P  pHp���-�����߀�� x8xD����_��~ "�G1�*�(T�x���<Tj�|�?4\&NAh��D�$�t���yx���|������U�������cjfnaiem���������=$4�GxD|BbRrJjZ����¢��_�u��M�-��}��C�#��3�s��K�ͭ�ݽ��ã˫�7�w����@����?���<"""�|����g "�Gd\1c�T���x�м�4j.�|�?�4ܛ�����_�����r���?|� �p�^@��3���Y�V z��G��O�9����>c,}�,v}!�����^���O����^���
l5Um/�*gFͮL$O%�ƈ�f�h2)�#9��B#��C� �B,���dl*���9�?���1rR�+�:������>�@��S�~T>�ӯ�{�}�9�;���H�e��S���>��
\ݯd-�<�@�zꏚ�]{��x�
?�g����g�K�W��>���^1rI���wi���Q�L�N,���S~�(_b6�f���?�k���MG�0wc8ń��ȩb|in�u��X��*^=2�vp�*B{�k�=/I�z�׬IB��2�f��t�������0����$�vl�v(�� ��|����Tf��C�\��#�}��S�|6�4!N�ġ���y�<.L�c��M��kW�����G�3���Շ 2A2�ٙ�pVo �
�y2���eJ�/2��a��q�x�RtT��'6m�gx"S�6̞Z���,��.k��b���m��t')7r��|/ip�Ɨ;��y�z�}��$Kw�_rE�-g� m�!M�t��v��a�RLv�@�¦L���q+���/L�l!��|턘	tEţ,�i�b�1�1�F��+L1EY�~�d.�n�/��G���|j�\�#8SK�Aj�S?���[�fݳ��x��r�Hx*��j@PӮ�U���I��TpYk�h���{�_�����Nr�Cc��a��n.��g!��������1���J��8k������c<�7�k��f��>�e���m[��RM׈̸&:bi�M]�޻�{R������=h��-��9��!�;���F���mw�Gf/ׂ&��lM�Z��az���"rVO������F��:q����Z(��t�=���KF^�y@�k����4��	��X��@�B�AA�dU'/����� 2ﾦ��h�8m����_��� �R=#D���kI[�|:<�VM��C�H�M�&-���ߝk��x�F�>�>Iq�m��ݦH_����P��͗�F}��]�$����aއ��-����-�gXR9]$����q�I�0!��p7\θ:ә;���uY��v��V&ؒJ<=�jV�����b7Iw�g�?���/5��
���re�(R�c,m�+��eX������a��!�H�y���ڡN��f�j��s:�����aX���H�	F���.բ�Ck0�,�̉��S>;ۇ�����5��y+�2u%a�%�lD���1��ދ�����̨�Mv6��(���ֶ?IK��iۓ�1����v�������
�OS�^��Uw�=ɫ�cĹfb�\�_Y�B6�hO4���i�@Qu����Aиn�8��2SR�b��Ah�T�����,�J� G���>4&�/_�?l{�N��u��sJa>+'S#
���56�@v�I�iq��ҩ�p�d�2��%��؎�f��QE�k\|O�H��Wr>YfӼ;�}� �S��j�}�{��ߓH���8��d/�l��+�	�b��B�_�nٷ�걼 ��G<T�wI��R��]�7��g��̈́ٽ��DG?�;FC�J�'Ӂ��7@�Pd'Y���R��:�Ll��kN	�8��?�6F����vąR�H�~�/S�b��]�74��ള&3D&|�]��n���dnWJ��^�!���3�Y�15e:^�/���!��_~�fn��|yG����NO7%=i�A�J�i~��Cn����߇���K���K�}g���/��(U�Y9�ݾ6���"]=miT�dA�c��Z�,�2-�Q����C�]����B#�:G�d�$+�Q
>�~�8fE��5�.1��D�Owkg�����6��>�f�*�F�6M���V#�E<k���[T���Uzײe�)B]����y�-M��M>����0M#�hO>�j]�bbO��6l�:ϰ�H\����j�1�V�R��������k�7�}����̟
������ɕ0q�}��*۵mg2��z|h��lu�m�.��.p�K'Eqڌv��m�W�+.(϶3�/�>.͹���N��F8M�/������P[=q�k�ʙZ�Eg����3m���Vm=ɿ�N]���]���}���y�b��kU{=�������J0����E��	=!!y*���(ђv�u����N����<z�Q�r�V�CP���8w|�=V��w��2�[l����Y�]��U�=����k�y�e>�ģ�� �}o�����b�����9����=��+Q쪒��Y���͏x��'��v���6w�k��'����8\��E�]��*!�����ڇ�K,{Ʌo ��"�p_
j*�/.Y��D���)�U�~5������[d�\�^�M�4!�6|^�1�9x�.uQ��� 9��nbۿ�6-}�z��H<7'q��NVx��B��{G���mG����JO������*��;�S&͎*��G.
uΚ�@����\z�)Wvϥ�:뱑8��äM�7�-})�|�f�R-PAW�y�#�n?�)6K�@�̩�9K^��p@-aGTb2�GH_N>kP�����Ed��3C�F��N�'QqeBv��dG��O�]&�hf��߭��uf��+�����e�ˠܥ�V���MYV�S��{����.�0�J�<V�v�ř��ŋ��E�+��#���SQ�se�a�a3e<������zt�D�����0t�h;�ڛ�����uhM�8Q�%]^�&`i��\�Ǎ^�h�o{�5���S� �ⴘ����ӓ�����De����Ñ�?�˛��:���W�ܻ"��0��V>�V�V_��(*_��<ý���[G#��q&�ZWk��!�\"2Mզ���@��ZB���m	�~��kKf).b�Q]�3�����N�1� 6J��B�M:m�K�^kv@)�����"�>�=׷6���^1���Y�D�KI�)ꩌ�c��I�֙� ��;!"�w:7�<ų��`W�YV=�w
�����������O��W���	�s�gC_ҥ��(�A���ː����;�U�?�\`S��YK�]g��*}зtbdU�E��12ۋ��7 K%��� C˿��,�B����E�m�H_�	o��Xj�e W���D���DY��\� }��H�]��L��>S/d8ކ�Җ�?���u�!��U���a3�St5�XpQ���3TB��!a��`E�"���Q�ܬ��9�4�
U�'i v���C{e�`�vV��̩!��=���?�E�=����)p$u;﯁?��cd�o���'��?	�[��i?��7�}UJsY���y#�Ҍ%ҿ\���{�3Q�&m֖<�K�kJ��cX)��v��d�+�i�!"�b2�YE#���2��Nijen4��J�[��2^*D��lˋ̶��dA\�9$�)Y.B����q��X#,'M����7V�;>��Y@?�j@W���Fk/���s�8���5��������0�uI�u��d�@�n�8Pt���ڃ�JѺ���~1��Wf�mؖ��M��߶�6��*0?���Z��B�Һ]�$[;���{t��8�"�"��n��}Jsgl��$@	�*�}7�[MR���3��e�&��,�"blPǮ���q�vU��R�?��cm���s�r�Mr�fJk�<��k��i�h�̂�+H �)�7�&��������4��&�)� ��Y^���=j�^f�%�T��^�|�}�Nܡ J��ϵh���w/	%Ø\��NCVD}~�t�yϝ��
�)��gz�$�?
b(�!�~���E���D�M9�1��1�r	Yg�ϭ�~������Ȼ�kV�zG{�3��e�(�R�q�5�f}��:��vB���G��R���QbhQx͟�G��ѷ�  �8�t�g������ѱ����
�b�\��Im�T�T �C�.�b�&�z�ࢲ�t��J'�Ǐ�J,��Uq��~�N6��D��j�~�9Z=�&�I��������9�|RHq�2&�B�7�(3HD��=~op�(�^ф!n��\���}bm�X�=��Wi��&n/n���pK��?B��5��/A�B����E�k�z[�\-^�ϋ��(�[�-@T��Ɂ��̖�U��4`N�w����<�-c�=CK����٠~yaH;�F�&U����ŋ`��2c\�?��M�t�Qi�IG�v�TT��`��m���o�$�b���1��F�P����$��k��%��,��;DpO
�[����Â�!Q����$���g�E�s�/q���h�`�a��T�o+u�W�w���?��L>����|јȧ�����J��	�
uU+\�&����6��<�*��|��̫I(y�������?��V��]�7�7�>��2.Ϥ����=ކ?{CǞ��#�>?�_�Ĵ�X��,�z\F�g�F5�2��O	�?A���j�����G�o�"��6ٖ�6�͍�<���p�����V&��e12+��!-i�QP�Z&�^�oR���P�Jd~�W�<\+��O��P7�e` �N����Z�X�O�����������V�(CS�0TR˄�{f2h9x`L�Ccm��)��������c[��lw(ʮ��T�=ɀ��٤�tXT�� ���3J#w��з��,��կ�u��ȟ�	���
w��
E�]8�%j�,�кĆD8������AC.!AT-��\*���)��y��J�ey6����gM,�ĐyĹ��
����}����2
��;�ma)�W_f'����w��.�I�ޅ� ��'�5����.e�y8���G&4̏�����h㷃���OgS�h�m�1g*X΍��|�<,uE�-|���=)�Z�Üi���d��`�>?��>> P�˪~Tcq�3�h��#V3qRW�lz�`����r��/Rw.<RFs���;�ND	�Y�[�:������Y���,c��F�3x�*��$@k��P�m���#oZȰ����S���T�[7��@]�!l4xoh�7[B��^� ޺�����Tj��Hx�yW&�>B}����LY�䍚m���]�!h�jȉd�I��l 7�#u�}���`��q�;Ye�JY+���
{]j��+[�2����d�w�7m"��:�#M#�\�'1��|���^�I�6��Џ|ެ��Hf�Ԫ��{%:�8hqxx��g��eu�x��)r���|��1��J�.D�#8��wf���	ӑ!�}���[�kt�f��t��J�8�w�A�hc.�L�h���?���N�Y��D&�}H�s��i�s�w��$+AC(Lx�:�P���'3Y Z�����Eh:2��~9I�Z&}4�م���}Yӟ�Q������"�~v�~Gjê�n�M��0Q1���&:[i�;�%ݨ�@o9Xw{G���i�s��6/)�������yju�Co6a�b='[�L�[v�+�h7�����l,��q��I$���O6l.c���~�I����K�Z����_���)�4�4n4O��V�O�#
�.���Xb'��ɑ�#Uf�<ɋ�-���W�L��������<9��:�)��e�[����B�]B]̑�4�%4Fh=#~��u҄��o��!t��
��,QFG�(��crr�|^}�1��1[ ��XL9;��t\�D�
�
�e�� .�,�$���GKNk�>S�*�H����(x�� ��x��GxB7��I+��}�=���]W�1��}���U~��Y�[���p����S�o��m,�G�)4������&'O��+L����f�B3R�A��W�p%��7����*Ũ9���dX���[{�
7����j�4Iд��E��ٶQW
v�oᳬ�X{�m=�7ڣE��[�ݟ�X���G�L����Jl�r�r��/wC��s�i;sJT���\�Y$VRi�(�Zgq�T�ͭb�,��k;�Z&�;��u�����R�n�`�-.�T���(l'��Z����T�,�U�7@�@	��B��c�e/�,<���HJ�>��A4nc�a!�Y�����@�Wa J�d�ˉ&��'�s�LV�\�!ËϷ�D�?,-��n2�X�rCI��4`�y�s��3R-3��
aQ�M��l�gE���#X���dB7���@�d�������U�M�E�ن�g��n x���#�P�xE�]覩t�2?sS�m��Sy�m�w 0�J{T�a�ZV�ML���m���KyU_�,CN��r!
r�`%��u@Va��0����x4B3���@ |��P`X��:��\|C��R�"��\z�""����3sx-����P,���D��P^�S
.c�Q"�\��}�׺��,�;���% XAkgs@��ܨ�H��!��J~�sɓ�P�X���YK��6񚝘6�@	b�@a�I��~�8j`��yb�Q�λ��3������Ex�ı��#���9�������+�K������,S���J���挒Ɔ� f����i���~��j��{��������ǛVT���F�af�MYe�b�����D�r��
4ac)ݼ�1i�'M�����",=#N�ԹD� ��ֳU,�p�$��]dE'���y+"�@���>N#�'?���r�٠���vYi��ؐ�|JӖ���pg�h�g�v��R�*Mmg�f�n�ڿ5*9e��
=�[&�\�ƕGO��~�@�t�?����y��7̻l+���ޘ|�̩՗tg��yK�ү��#�<{�ӑs��'�8C��X�����Aʉ� .¡˴J'A������;��1���(�)\�j�W��#��u�_n��TAL�Z#�������p����q�!��3n������zڻM' a6��k7�[V(���Y�%�0�蛣�2Ee�3���9ȏ䀺c��Nsj>&Пqy��֌�X	F�T��YO$�B�(y�?����Y�����+��`�Igs�<�;A�eS�4���p!��.~F�F�p@��˴�����z��g(�ۍݰ�I��ɴ="�*a���VkM�Q�AUQ�\����|爞�w�n`n[&��� 4�;~�%e�����V"��mB�.]�)��E�".C�0=�eJDj]޽*�"�L��
~8՗A����Chd���j�����H�KGz�&�49/�CMT�;��L��R���h~�o��Q&�N�\����M�P��(�����w�L�6�%[V�.��d��9o7��H�ѽ"yl��������/��#�ۼx���W�Ă�4��ĸd�HHi��p혹p��i� ����Q]�dOK������].E�tD�dӯ�}�0�Ć�,5^�Bh�A#>�2�QI�!��Sؕt���]$�?f��5�	�<^u���団�k%��@�������_���5�a۪i�0��&�oj{�OzG\z��T�(���(�o�`x��s�p�U��i����i6r��W	!��j�:oNh׃��f��zh�$1����K�1�� |N��Z��g�U�^��˽���ڥO�lm򂶟���]��c4_�*���(C�6��RX50�Ό>S�F㖒�շ�a����m��RmuFe ⧎	��[����e�\��a��u͜#��:#1E=���N6��������`�
�&���.��ЪX��MfDwM�|At?����5a�A�S_��~Ǣ���^�t�z��!�Qߣ��Ո.gL|�5����b#�2��~���xw�v�)t�'L��B�Z19zQq\���-&�n��g��R�e�i���b(��s�����q�wL�+��{���u��egWCc�	"���ϗ-r�ĨJup���c,�+�%3� ų<5�����o2���S��W(�)�S�g]���@�O:im��5�.^fg��m#�Ը�Z).�hr�äh$���t���X6�[�cـ�6��c�B��$
M#�������2�b�b7��G�һWS��-1�ޚ)@f�I�g�^O6)��|�SxT�ۥu��<�����'aF5��%�����휩��� �x@���U��R��T�p:�J�������T���du!��at�)�ҏ�k?��F;I1�6�m���GI	n���r��;���0�`���q�b���$ܰY���-_k`.����koܷp�D��VgM+�pP�,�`�*�J�{W��/-�SQl�J00�yJ���f��Ƌ���d"�-0^�72W�<��D�NR�s�t|#�������̤�4��uĥ�kW��D�D��{�~�9H+�0o{,�)����S�~	X��*�NfWP 8K��{�G7� ����v��r�W�3Vւ�0��bW}����i	�n_�Z�ρ��W;&6{e�E�CW���
�*�����K8�P}�ǧc����X�8�,R�����|��y�Y��rr8����?�'�R��kم͸d${`��BF-;�ؕy��L>�+��D��J��1v�Oа��kv�����-F�@���/�
�_�q�M�B�h��M_G���Y;�|����Tq%!��^��Snj+�]n��y�~ �cq�_�ZѶ@�r�I��2H*���)��7'��w���x�0�'�R�a�9�}���H6(���)�oq�T�K+�$��Sd/���]�,l��7@�O���Xq��P�iw5��%4c��d�[Gڹ�z�p٬�wVVw�z���e*��J�a���a6g٤�I K�#��w��D����p���Y�=^�!;ؗTb����`+ئP4��+�ajL�a2t[�q�tC�΁��?:� �7QP�Mqx��|̨X�'ʼD�ȧ��r?���33%Z���l��bLTox��h;P�8��<י���ȟ�J�Е*QحW坕��w`��ԗ@�����o�[7�ߤ^�Fsk�k��� l����@*�WШV�h�!���A%��I�&$�{�J���v������<V�ҿ�����ܑ�h��#+ۣ�-iܭѥ���KQ�yF��'���i��=����&����݂����j��C�S�F�G�z
�&�M��y�,�V�f�`V���>*}��H=V^�G�m�kw��3�����DM��#J�=C�!����\ c*
���}`*�X���29P	_KgU�$-u����@%��  @%0�ր,{��K,zbw�n�q��L|��� i}��a:��s	��8�U=G�����FYOg��&�=�k��$��+R�X�Y"�]U
k�84�����]C�=.~q�z�9IGG�\�*��$rP���k���{�����3r���O�3�o����`M�oU��V�ۃV��y��E��f��{�x��;�w��P'2P&2��������pm��i�Ӈ���Β��&)��S֛��>w<����;\���1���k/3¼����$b���b����ap�J+ލ��̇g+��I^����V �h�DY@�%Y�sR�P�H��?��D���`u�m.�Ȑ�B\Ʋ���!@�&H=<zZl�I��P%nq0�}a��p�V�����R&��	5�-w��T�[�����TXL�6�mƱ��q��m�[<��t����7'@� �AK��T��l}F�ߕ�ӭ��n��e'�F��r���&�ĮX��t�`z�mTB�Gm��H51���*J��7������=�TW�L7ɯ��
�*،03VT��x�j�cr��� o��F��ϟӆ����px����6}l3��<�gf�9/���:n��)[�����q2�J:���jl܎��!�z��c��U�m}^ݪ���1���\j��$��m8:M�  O���uR�
]F��>L�b��fF�n��kɘ���'z$,��ՓϿ�A��2�ki��v�a��<�gܤ�U�胏��S�%��'��3���ʢwo������|
H�˶�W�{���_:�jҮ˘㗞OJ�ƙ2K����1�#K��%��u>l��b��.ּ�W�?��:���s ����2(���5��U�M��{�3�H���+�!~��l�ɫmz�|2��5��V���& �E#`Sfr)�A)Y��avp(@�c�������L	�5�e�1yN�A�HG(� W@�M��l�^Q09�2���7Ӎd03�(2s��g`���m��0�T�շ[Ep�Pt����.U�pʡj!��k䁙�L�3��#M�B�$�cn�#�J2]ܔ����d��,'l���S8N�wm(ug��3��Ͳ��4:�
	EW��|F���]p%Ĭ��*s��+&�^YxI�7_5���~-��yuC��ƨ�Vv<�(�6����o�6׃���:3�&��+W�|-�1 �E��W��w�~��U�`kte�{g�m��V���foNPJ���Y�/䙉T�6(P�)bU^�Ӹ3 �x�����}x�5���������d`d	ww���oڰޅ�b(L�������MA����c���͎�6�*C���Ǳ@^�$^��3��,	�$��*l���8�Y��)Z9r��I�E��*�����}.�"����ٚ�޲�����%��J��xOP��} ���\�~�(
�rF)>�-?h��0�BPX�9���\;�|�W��9?(-��q<(��,�E��ٺ��I_�l.%��ޣ�����O~�p'�h] ?�1 �O���+�h=*�ÙseL޲$Tя����T��b��f��҃<tU�t�DT
�(�c�|
��G���-�A��G_���2�Tz8]˴�~��
/t��sE��<ت�	��Kd!�`f�%al��⩛_4<�Eu}��RI���Q��[��#�2�`<Sa�4W���?��r�9��Q�?��~U�M?�Yp1�)��G�ּ�5�=e]���@�Ҡ�� X"���z=IHK?;pR������9,�vd�A��t��ء�	�<����&�88�����/�-f4�*�1�䆟k^2Jơz�!���JI��K3��� ���.o F��;�N�a��Oa�BX����e��)�ЍR.� ";��!:���_���j��� �F�B{tYO]W�:Z��zr	�Y[m�D��E]m�y0�v'��e��I��_j:�^�P�֮﮼��T�24�^�̎Ԁ�����`�j�!�{��ʼ�U�B�>�֮��]�i��&y$�� ��_��Qd%�6)af-j�j��g{��@>dYZ��	N����T�F ��!G��j�r�H���2^q�YO���u�3lĊb�����m�'�+(���#KҬʪ���mdFhS������s�C!�`��mwh�L%����:����@�ƃ��t�t����֊q,�nm7|��$���>�����i۳��2����P�0_�SeƏ����:)��1�*�d~٬��~�֙QS������R�b����B�ǽ��D�I��P����*�T�0v 5���F�Mq��1�G��j[k!/R'����#x�h�#��ͧ>��$zl4F���d0�b��鸓��4I"���V.ؚ���R|�H����p�M�	�iAL�i�����ڶ�q27�_2F�1 ��j�e��ZN��nsNn�>���NmLܴjl�V$����Ҋ��e��'u1�PW��kcO�7_�d/�b�m+�U�ËV)-f�P���r(Z1��e ����S�zG����s�8�C�񃖺��@��� �x���U$��$<2˘`LA���T���CW��)K���^��N�����D>���5�s�;~{�wPb�4�*��d���b�I�9y��bmR��4)"x�[b�qp�9 �:*D�&��Q��m��&\ن��!���ZR:�˲4�ԑ��0�U(; �9jT�e�:��c7�`o�,�����YnCn+�Q��־��t`�;��Ԝ	�&OWն;��h0{��Z= �S�
6&��>�	�b��+X�r|l�R��ɋ��8NԜ�I�R�?Et�c�yx;�����Y���n T}�I�y$gjp%��B����WL�bD|����N�}����Qü�o�oV/�;����|�m�
9�M	{!��n���ڢ ����|+s������	��EL%,�:eB�;���� ��� ��<h$!��l��#���y�2ֈ�e4G/����s�N��#M\�֛;�(�W����^m��]�>�7���f-�K�,%��!#�lʻ�`��4v����������kBR��=j�,���2���m�s�h��B��ß[M�u*}���R���B���)���ьa˷K����~��馌�.{����R\}��(b���9n��y!�2�����Ͷ �ܔtҔpdٔ��e�>t�[�*bX������W�O�_�rE�=��3Ξɕ��#j C�B6ս��m�Qc���m	���H��g��)fIb>�B��J62�@�9�uh�Q+��4si��c�=�
�l\�Y2�'�i�@��)�L�Rmn��@�^�`>���u㾀q�ֲ"��_��7����i�S�ቂ��¶���q�ЮL���Exs�X�W�&�vS�[Ä��K,ѡ��EE�-~gq*�e�H@�#=��FE��o�}�̷%��*㿉7g�C�Z�<��&eC�(�BO��.��ZHlcY�/��H���icNIU@�!������U�P�i��%2�<���P��l(���=�Lun�i`?mh�S>֢4���!޾�kn�4�Yz|)3���N�0<��d��� ;ZIH�I�"맏Ќ���`Q��L�[4�*�sl<(�v���_
�Ǝ��8����/$A��oƐ�q�&�	0��Ax�$�j��T�zf.hib����!�(�� m�Ϙ�1EA�R��_��PL����cӡ�Z*W�O�����4���)�ʛ]�c��'.e�6οϿ���+��ɷߝ�z��r��i�q��;5.��TE|z|�9/l�S C���ϵ"�Q�3��W�NE�z-���e��8RUǎ
��.�VAhNC�HI�NFd�*� �g�x�d�ч�ςZW��%�B����E�j±�3W�(���zm��>x#�n�_g�N��1N�j{t��~�&V�64c춀�+��`�3�7�S.�Wz?\�t
�kUv�5�s������������23�E���噢�X�ad	��)�%��j���N�]�ٴ�u���Q�o�7�wɐ�ͅ{��98O����;�a7� a��d��i`n�Ð���]&�8:��^v=�$�E�eM�7�Q�Gٷ��4����`��m_���܆G�c�L��{�r�����Ĵ˾�
����x>_A�>9��`i�x���!�z�y�a&�;M#���+���� ����S�S^6��}|���1��΢,�o�����(�1�LZ�l�ƺO�fT����U���qq}x��&aBϱ�/�3� �.�X���U�6&�p�P�9��ZT��8@��c�a���YH���@�I�!�y�ڵԺ���ʆu�~��2�*� ��H�]ՕFӯ�V�V-0�(azL+����%��q!A>����2F��5<���&���m��q6���3o��^�8�C����;x6�>(H(@L7�����ʖ���_#�m��̨q�C����11�컑y����A�S��c̈�佇�g��%k*����e�����%;�:0u~���l��h��v�26����^��ƅ���c$�.��Xv8�4 ��7F^?��3���Gg��������E�򭯸Ga@�  �当SU����-δ���m>�/2&����I~��� ��T �k�uD����[�+��!\�R~O��6�/M��������Nf�L���9"�������*�9~#��(ʩf�UA�{�9�I��i �S��z�9� ~��%WP���fas�I�Ѳ0nQia�Z7YM��K�'m�Þ��
�֕l`��O��z:�/���B	��AG���՟6�l�ڍ�r��r�@�^�&s�2=��0�d��mp�&v9����`ږB����c�S�W��PfM3N#�� xiN,=H�2�5��`��;�K��ZV��qulF��_d�)-�Zc4}	q�I<%}�n�-`���Xi0p����.4h�4�usG�3Ʒ� ��x9���a}g�(�Ir5�m71�Ү�0��W2��߮Xػ]�Ge%,�
�rfO��ԘtM"����Z�F��M�6�K���{]=�lH7��Hjx�q�nq���O��[a�t6&��B���tT��e���ߛ���}���9��-_�� �n Ͽ�pz5ןP�P�@�+���R�C{�._�����n�3�u|o+��9�ˮ�IVǎ�2��&�}t�i���ػ��<J�����N�h�T�{�����M��F,5�G!� !��6Jю<��m��ݳm~Će�F�c�0vtFD�i�J�ԗ����.�ib�fN�#_j�eƞ�]z�hί!\L����7]P=+�R�9Q#�Q#�0Fw`n5�����H�����l���ծ���/u�=>��D'*B2M4��n��H�D����,tG�9�g�l/c��\����4�Rc?F64��I�::z}�+�p�r�@pD�Gge��`�I��:��bT/�]Ǜ�0�$xDO�r#�ek����Eb����TTp:��"Qp���`e�FI��Z��fո]W��(���;��Nr�늤;�1bN���s�=(l�PgL�d�";�
z46�)����q]'�~k�/@�d� 0�e������a(����[f����l�5��1/g��Ƒb�*^E˖$�֋��m���m�Ǌ�H�5߱�S�����4@���9��k� RQ�&Pwl����d�`�/9�ޮp��?F�A���"�Q�P�ׁcy�+�L9L�m3'X��<��/7n���]ӱ3�_���,l
屘;I�������፷ld��#k1��
��0��PѴcaQ�En��Em��V�#թ}���*�UZ�dX�"]�]�쾽�r+5�����Tt��I�Y����X�A�-�/��	�M˕!.�c���v#�����1�4p�F��K*U���)���rƒX�Y1�&��I�ݒ��x!���Et�{��%n�4��9����C0�I�G�f#Q��E͇@G�2�/ZIg�/���1�K⥴�6� ��_�+��A'%n���,{�~V�mm��G:{� �v �x�d�-	3��c��mt8�=o��Nۘ&b�X����6�����-�{��<j��.%�~>M��v�9-�LDE�!Ę���]F����C�!vMX�%�N�&�K����$��T� �\�H��taag������)��F=*�6"�<������lr
�}:?;ʛ4Rnc�X�ƱP�0��y3�%k~{�O�O��$n�7�Z���X�aQ�)6h�i��s����ۦɘ��!����s��|$��y���Y§���r���x�A-��P�Kx#���co v�&k���L��+`I�(n!Ӹ���͠��W�Α|�f�Nb =\�L������_n������7�Tu���:���ZW�A
�sh�� ED�!�w�iW��`)��r\U�3��7 *���L\.M��h�n¶��y�Aݱ��i��A�Jvg�GH>�M��S���K�E��ڐ����&�;�X��~��v�Q7�#0����p�e�@���0L��9�#�rW�̧���n�k���-�%�����l�!N��H�ڟ�̔���l� ��_�,�e�?x&���%�p���v��H��������]_+��u���cxP�����  v�O}���^6���\�g�8���M�1�AQ�L="VS0΅͎�t�HG��pz=�r����o��CqE�a���۸�?����qwrj�6��]�5��'�!ᤇ�-C<�*WGO�|��E���A�qOXp�H����=O��&�[��*��X�� KL��ϒ��4���u�VAq8q�� A�� 	��A�Cp��6�	N�wwww0@p���/[�Wu�w��y����JU��zR_���n-���a9��7:j��,K�:f@U�X��]{��{��ܭQ���
����y�(䮖ޱ�-i��O�7]���塰1��[J��\\�`l��O�i�P��A.����ܒ����AM炞���*C��p���D�l�Jj�w�~�D��̙x�
�9��f9N�Iψ�	��#�,�-�nk:�!_�%s�6�J��%JZ�g[Yy�O���������]���7�>;�@~��͍^�-�!*�d�N�f�LȱӦ1��k����ŮTR���������+���B�s�5�+�d�8nڹ�����@�����?��p��Yu��vx�.���vձع)�s�]ce�B6�QX�G��WVyB"�E��b8s���\�蜇|3̎�7����䞌���%kt�O2@�>|���҃�`�����Z�;N�1^��+��v8����m�X�+e�"ׁ��B����W��c:��s��~�7�'=QӼ3NU��C�X>�!}����m�O��`�M�B%������N;��Q�cOw�M ��ׯ�$�E1����P햞M�j���5����8]�Uy�CX���|�9�� 2�����F}����m3��7}�E
�
~
�.�} G0ʇ,��D�C�?kE*��A��U<��PZ��w��XCR�[_�oW�+�<D������fv����z���6�����H^�ё��U�i�!�e��;��f�g��q�޷�K��~>|�a���DT�K�s���݆L2�+���~��47����͔Ckx�Ge%����l�>�6��2���g3�_��L�ς�o!
��{���8�/�њ�0��c�ݎ�`��c/���%�柙�8�J��Zp�or�Q��x̹	=�bd��cm�g��!��	�C�7iR�W2��l�M=O��6
�?�*����J�Z��#�L�������>��#�����O
�6�C��F�Հ�s8rm"��
wsj�fڴ�)���oOZ��S��j�6����[7�ܨ�]&�7!T��7N�I�b�qw9������c?!َ�y�E�K�$뫻�D�g�������b�����f�Nm_�r�0����i�~�h-������ʏ����u�疛2۶S��rX�2��m95�j�K�
cK����=��h�eʛ�)���ˢ��wp:9���d����en�� 3m���Ճ��랯 LV��L�ިr�q'�Ƈ�R�$���/Cڔ��-����߼����(����/�y�zԇֺ��ۏ�ˣ�J?��@�H���3q�v�Bc��)��Oʹ�=-7=�ǫޱ��$�V�KT'%_ʞ#��T��,�%�z$S�Z����y8��}���]U͑1F#�<G�w���[�!Kx���^l�Q\���L���W@c] �!������@�#`bF��!��YeF�-���<��:��`�mm�n�3���]4[��Ǵ�� �	-T�� E��,ߣ4�AC3%4����s����w���-�}�!�!4�os�,i�4�W�'���<m}��S�-��ʦ�5{b���v��_N��4�#�FGͅ�w��p`L�M�e�[�a�ڽ�4���;��*���[{��z�ж���k	���j5l'}U�5,��|@��������`[���P��1��n���UZ�8��7$*/���[��y_�bC��0L`n�N;�|8.gb�X+;�n����s�Fwi�8�����`����5VE�I�?@ܹDk�вh�ޤ+�`O?w^���n=B�b���w>�`4�5�����V
#��p��1`�qͻ�и�o3�i�,:dݥo{���\�4_���k�:�+�o�\0��	{�	0���K[��~�v4���������1�����6.ܣܻ��G9�iG�_�m���+�T������܅A_'&���m���m���T^k9���t�j���єC��9c���Ƹ���B��cp��"!�`��}�H$���}D��˫��%��G{������b�b'�J�
�چ�C�])�O+��n�� ��u���`�X��Q�1�VdnNR��AC�/mm�W=ܞ,�4���)5ĉF�I��i/���
0 �4��6��Hs���ώ��fN���s.,��<N��md�i�ƹ��(��k�mȟo5�I�M2M*U��ll����"*�D�]0#����IXNU)���q�>����?��t�%���-�IR��)�퐑=�O̶f�J���HJ������$X?;/6�r��
(�웾ڲ�i:m�Q*0�c�({��(�{���շk�0`��B{m��`(_��M��c�Ob�x�Z�
4�GB���w�e/�ԟ^�fW�ڈF�v�D81]��[�p�}t���jt���6E5oR�K�>�Έ�4�}�(ыP��8�Uԡ g���%�� (5mc���l]>��l�Pf?�U�R(���K�CB��nNF��d�K�h�D����J��gꦟ��U����0g�i�Ge�A$���̰�A�Z�c����z�+^#�I����g�eaE�^T�z|9	tS�����u�S|��s��-�z'�WkD���2�n
t^w�/�׿ES��W�=�,�-�+�v}�U�N.o2�`tSPm���8�[�fM4|� k��׫�e�B���\Kn�0�X����w�SYQQY/���=1}:����(�|͘i?�f�|Xgx(��<�&Bv�f�䙴k�h��s2�̵c����y$y���'įΓ�TP�"�Y��v���q��k0R�Gjv�9�"B�"'W�K��)�и�L�W�����^"�����D��T�,�4Am5�;k��'}2|#��K�s��R����9�&b��}�4>!��n�L⹵sq�}�Ye9�.��O��C}n�7�@M��U�>m+Q��2wY��4aS&�!�:n
v�>'�N�M�vch��S�I��S3��u^�E�U?N&(pzN*	�;��3W:�_y4��Oݕ�8þԡ^���|�����
�b3���o��4D\���g��N���O�~2H�ܑr��D��a�����v�|�@,k1kAM9��h=�Ƨ���z���6�ފ^��̹f��$E}ֺ�mf��Ƞ��.}M�,�u��.�+����Ǜ����q�G���'��8�L�� ��%�'��fv��d�+��!�:���,�L,鿩�����^�<?7�����Z�R� +�����d���{�ϖ
u)��ю�4M>��~O��UJ0��$Zɵ�P7��wWv&�� �[��1�}E�;s}�xL^l#�3�+��Bl�o�b�P�Țh�K)Zo}�g�T�������%w�k^��:�<*���؀'������:)s� u��H\A�-%����dC��3�J�86�KDb9tT�.s�`�/,։�h��w����4	�]k�y��.����֚���o+�؜��\��k��n���V���Ӭ_+#���W��,'ߑ`.��^����U(�챂D�1�qy���K�e�D��#��B�,'I��W}(�,�,f�<=�/�0����|��;M��$����]��([4fڈ��ӟ��o�gG�ʦ��k
��7��5�,Z��&�(��3��Jh��Ժ�JP���MR���H88{��K�-]@���;`����o#�w� Z����X��p�	�ל�t[8l�>����9��a����d�{{���c���G��	[h{�Y��'6 .�jPL�p�����~N~!�/H" ҵ�5�m���l��P�̅����#��B�l�t����a����7���܇-2(F�;%{:%eKy�h�z$(�g?�t6O|4Ώ)ʖk�IF[OD�F�y�a�.�*�+�3�*w��Zw�[8_/I�DGF�d#A�eD`Z���Va����;Eǝ���V)���\�+m%+���8�U(.qx� �K�d�EOI������R`!�բ��Tq<H�0L-ԗ�d�c�<��+@ƒ19����9�V�>��z�ܧ���"�l��Ah"���(.f!�H��� ����%�=������*CJN��gv�Z:F7~v%d�����}��~~m�1�Ʊ�)�R�S"A���4)�O�/�q4��g�w�cӲ�U�bŊ��Ⱥu|����4E�b���R$AdKÓ��]�-j+����;���u���4,H�X~A�3]��)���ۯ|��X�y+ �^jք��L<�#�i��M���$1RX_&�_�����P,-����Q���|��w�F��'�+�K+�#D�Yk9i��d�,�'囂����'�9���ߕ����^L��/���.h�g�W�0��+��0�llNT-4����}��1��X�4L̽�/Fe��?]���jz�L~C�Dӏ����L��e��<9���f�:���/�W�I��`%�j�9C��3��.u]~x��/B}P�9h�#�K)R�<ɬ6����g��N�W^��W�U��5ҩ��a ���,���Lf'XI��]�"*�÷����o���������51��;g7��9L���@����0� d�@�������8������䲮��;�
8��N�!ڢ��M��#�rM�_g>-i�a��Q���M��W�q.���D{���E�5w|{�����#ѷ�S��ƕќ�2���F{�K�-{�4���R��� ��M�+�	������ۅL`HJwd���W�&Ns�0��֊̨��6>2�����}X}F�x���`�5�s�Ǝ�"s����߱��CЪI�̌Ɛ'��a��'~}C؎"o[ډ5�bd�=�c$Z��]�˂x9.�~Op�flt�>g�b��n"���K�>1>��!Y�N��^���T�B/��ߑu\b��0V
'��\�J.g����u'�#"���/�h3*�D�֮'HݶnagɷO��v��~��K���J�\q�:V�5Do7ޟGRU����&�t�x�y�)]�7C��[���b��;��Pu�U�>�cy=�X48��n�Nߜ�s���.����_�'?�F�	'���t�Q�_V����A���:�?�*dOmV�n�T$ f�K�$it!����T�(v>pg�h3��wg��� �w��h��1Ⱥ+�i���CĈ�1r�@�Z���lp�B�ͮ�C/�Q&���;9D���%��?%����O��ߕhb��@��eiA�AN���)��B���5���gu��%�������%%�!@#I��J�t_�(���~u�� F�jb��:M�l������G)�%�TEZ����,��\�hts�ڎ�
�z	]�d"�^��rB�u�q��w[�1�*��.y��n ��:.^!���g��b�L#Y��֓����ã��5�$*��_У��������zx���\���>O=��!d0[pkdХLG��_��}�2��$�q�c��;��z �����ᨵ�㦮#<w�L���`��曩%������FsZйrq��T[m��8�m5�2aa0N������8�/�a���)��m�CY�U�\~�׶�ӑVv�������D_���s��ƪ�72�o���P&	��7_��]��*����n��f���E<��,k'���v�{����Q�CJ�D�.-w��
�ۖ�nm�w*����X&_����\�%"zjF-�`O�@�݈�!��k�s�]��gLu�Y�,��6Rlo�l3���%�����䍝и@Ffq��āSύq�>a����P5��<#l�Y��Ç��:�ɿ��o8�� B��lxp+�T�M]>Az�Q2mG�3仹���U%���4���X�[ڂ0�c�����Sp��G�����_��
�z�zn0�K�2`����B7@�;d�du�0d�� ��xqò��Tܒ5&JXa.K�mH�'G���齐�����~o��)��E;~h�ę/~gM������P_�
[?a+�|Q��������ިE[�c��m��N��S�d�
 ��C���%+�)Y
e�v�m�ɑ�w�T 8f���_�Z�bϳ��,ߺ_���Һ��U�҆;
�eFL�6M��?_&w{�A�CR����� ʉ3":��x
��L��2i�6Y:�����m��ޠ w����n�pIq�^��\�n>��׷�m-�c�llTln}4�����4�K� �p�Fu��)f�Dh��)�\�KI�8@��a�QR�e(b{;��ߒ7����$|*��jXBN��&F����I��2�z!�ϟ����J>���l>U��k��gAX��D�����I��-lR[ʾc���IX���7�L�^��7�/�U�5��.0�nS���[rMI�Q���Y�1��������ii�}��3e����u��
�2�,�di|&�n�8���FzO����Ȧ6��j�).�Ϊ�A�(W���}���|����xF��h�.�u�%��b)����C6��!�u�����U�����(�Vow	^�i�G�&E��z���{A`��W0���s��V�9�Ȅ�۾U7~�O>E9����ȌR,� ����΀eB�ɑQ%�%���m��yp���\�c�:�K:��
�Rp�I��L�"<*=Ҿ�F��mM��w&�����;glc��)�/�m��r�z0֭W�-9���Ӗ�)]�bb��-�NaUn}�J`�A��+}���bL�ߡ�I�ˍ/阓��q��7Ըσ�����1e5�3��9gkh�>G�
o5��Q��ω!�I��g��)��������ri�6��n���Q}�|��	��-�Ng���|�a�t��4�ȝ��������K���¯�Ԑ���w��;s�nZ�OU-Ћ��Ѳu�����RZ���\��<�h�=�@�t׀��-���,c����A���"Zp�w�Rf���8PoW"#�,9ޡZ�`���tO�72<��6&Jc������o��E|��5�����KA��@Z�ł�g���qK�e��Il�ݞ�u�cN,�~*lE����0̵�'�����U^���?�G �l���k�gj�Z{�GV��3�A+2�=7�,ߩh#��7|W�zÀ��JH�x�m�,��w�i�o��~7%�sK,t#�L{�MEg!|C5	�`%<�|rI�5����i��E�6,�_;3f��'�	����b%]�७������sz&+�S� �g`8��]z:#��uNE{*���"Da�k����c��򧛑� �(8�Q���i�F�UU@�7�u#�����,�Q;u�B�E ���7Dp�����=��t�p����O��6H��1�c���.�^�����!>����	{�ח3�����OIY<RbG���<�R\P��&���A|ŭI�����_�&]ޒ���j�W�r-�wѧǑ=��0ơ��0��U��+���z��k���/�\��U�)eļ����e�
uP(��7�-�!!�Ve�<���˨xm��P�C}�����ʝ�@���)3|.�iP�v"�NGPR�H���7��d�'k��
ٱ�u`��`������L��ƌ�;N��r��<�{>����>�
J�H�O�kq��i�9���A�J)�AFm��1 I�/1n�]��i�~�9�qr�1X��>9���6!��ȝ/��Rʗd,�m���P��$��w�[�O�~B��x r^J��B��\2q�ZX�B��;1l��O�G���i��)��P�T,����'i����~�}s2�p��%���heHC>od#H�|�&�Rp���Ȧ�~U�L*`z,�Qn��)FyΞ�q����9�3��ԁ��Gub�$�p�cQ���s9�q���,yϢޤV�2��d�mP5^�p�Y���L�
] �����Ɖ(z�_!!�&��^(>�V/1���\������MELwE��l����G(�JA��z����\������/��7	������6��$���?d�b���r^H@����;��Uz��L��P?�G�'B�6�??y�����0�y�-�Ꮵ|�tL+4�k]ƍ�?S��޹��� k��c�I��K%Y9[�/�%P��n���ſ�<�}�76�җ>�NPd�T�/�sld���T�ẴvFV���)y���a8�\�ϿP%�,:l��]���	3���[����!��ce�_)pxs�Vc�e^��K�w��p�U������®��?ʹv�`.b����MX���;�� \L�ێ,i��_忓�s{�j���_�Ô|NM�!D4J�+����z�7{3-៩z�l����y��H�jH�1x)Ͳ����̆�xa���N�ef[�P_��go�!#ղ� �Ok2S�(��<�D��0��H����휭]G��II��)����U[��?�:9�ڗ���������ۊ�G:�E�de>�B���Aչ
BS	4�Ұ��-/']�_��[*���K���_:���q-�t���Gz�ņI��jl-��	����[�wx�bO??��1�q����Az�S��o�q��p����b�5��-I�n����D��W�;�y"�y<֮~1��f2[pޔ����x@��	���w�m�'�!�[Z�b/���b���n'4r$���h���e�WG敜����y1g��#����h6�EL$p�Q�bڄ��@N�蟛�e˷! �M��ܵ��ܵF~�(��]@ �oD�G��=�M��&Wa n\�k�d�/���\��L��DK�z�E`�2����r��	t�M�%Xr�킞���UGp4l(v>	K/����*�it��v�z��fu��;4�SV&7��6�<E�P��w���%�%:�ܧՍ\��@��-ڰ��zPT�g����cr�g�`����=�=�	~��E`������P���8S�&�k��>MA\D�6�>��4'9j�,Թ:gJI�*"I�����d�������-8� ��ѓ�1�Py������e�@�D��q��jL���Gq��J��>�u����Z9O�{�i�p��b��_� �8z?��x���0��P�j��2���Dڧ�j�s��� �5{r^+}��jM9���3E&��%��7z~XL;���.���z�^΃�}&���ey�?ئ�1�T0s��q�K�L�?0�]Y�a���?��������/�}���Pr�A"9+}�jC�oꛝgp���� ��`��n��	�Լ2�:����}�;+��s��������@N���m8�|b�w��O�b������ӗ��-��G�� d,(H��>��۠�s�����F���3ts2� �0�ܠ���-�U�O���XO�s~9$E�����Bw(��X�h)}_x����녓�&g��26s¸�T�n��4/<:fb8#����4V��l) E��%P ���"����O�5�%����o|�G��:�a��!;���%c?�����结G|H�F��W~���ey.}B��b�X��Y�@�b(�s��¶Z�%�M�٩W���4����P��Ri_tgl�����I��[��\������d0��MZi1R+������fi����<Y<�=i!R4|D��m�'��� �T�3\�٨('G�ܤLc��-�?DLϑ{ϣ�<��^Vf|� �bQ"¹G�ũ�s��f[aq}X�Ŏ��,��R 6�%�K�V�ఠ ͻ�LL���B�w��mQ�����B�j?ȼK(xN��b�k5d��'>I4���d�Wq�W��wV�Y��3�:�KD�0H��*Paw i�C��Q8&���>,sX'+�%P�~2��JZ�F��=0F�Kʁ�Σr����s�U�]�+rTqӼ^�M�TԲ�I��T��5=21O�o���Č�{�M<���DS�hq�Ƒ�������<J�����?�M���9òeۉ!w���N^sW8q|�ɂ�;�"w!�5��\��eW��e�Q6��S���Q�Ta̘�H�L}������6$���qǻ+���X�*3�Ckyܙ(h�����1���B��r���/��Z �!����c�ּ>�n�u�<�v��<O�c����I}�i>�;��l>�d�!���dF)��O2�k�^��֞кH[��7J�~�!䷷G\�ċ�N:�^���S���fMÞc���o�Y]�T�m��Z����TÑ�Є���զv�Σ�c�Er�N��뷘���fr�TS��D�+�7/G��Ѩ�]ؘ����j4��~�t��V���Qv]�Z$O4ngR���)�ŕ���Bf���.���T/���+`&
dT� �����v�p2���L�����k���]��#��Om���[�t��-����B6⥹b����$Q$]�����8Ke5�V����yޡ����Bu����+�@��ґ�6��hd��+��.�NNyw!h�<�;]�e��V.�k?�ծvp9s�?
z'f�R
�>A�drM���0��$���Y�Ѩ�D⏦h�KԢ�/8�Ʋ�@�b��;yq&�u��ҡ���+ ۪>�$	��w��,o5��<z�Ձ�^VB�}I�=��Čy�s�@3��괐�ːZ~�,_cd%��i����,e�=xt��N�K����T5�sԻ�-�]4��JHB ?�E��r���rPM���[��n���{SaӤ�)T�o���rl��t,����l��$$3��=�q�j�������jO,�������Um&���ޝ5���V�{	t`ХJ�y	$�0a@�>�������H��(�]+6Nq�,W�'���q���Rا� ^�{P5J(]݅���V��� ]���jw�}��$�d�.���]��F/F�&-B7V*d.�iP�k~��|���r�:Rۧ>~�����ԍ֫��C�=��/՞��	,o�&�]����1���� t-<t��"�#��D�b�a�������oY�[S����/o�7��MD[V�^,ّ8/m5����E����ܥm��ۖɹ�A�B�oN^K��O��P\�z�c=��Af�Tk�~R�5�"Av���;U�O%�\M�`?�	��R�Z��"�L������u�b�n[�f�w�����fG�M��(?x&�9S����p��V��KH��kN.�Q���k��qQY�����ψP4��$q�ġ�l��h���z:X��2�8d̂`�L�O.�wkcIZ>����Wm��I�(t�^�M]q���t�Qc~x���լc���w��d�'͐�5W�%��7N>k����l�����q#ǌ��^Mn����=��HYIR�(/��$����g�Kv-�����(����Z�uAЮ����t�`rZ��z��APr��;�|����%�� �<G��=��Ì���G%tM��?n���Ao�b;�c�)�-��������/�m���s��;�2��P(�{�
0��F�� \�2fF`KV��n0w%��� Z���(��@��xI��#9�k0|��+`V�4�VYqN:5̖@?G�XS X�J��=H7	t+nF+���^�(t��x��࿉u
t�t1b.�>5���/0��ي�;�����ej**�a����7a8�x��m��V���h��l<Vĝ�����|��0�ݽB�y(#8@k��;�"\���$ ���h2�B�i�B����|g?������i�ić��ns���������	w��K�g���WU��t�64��S�]y��쟮�
��f�����=]"#��d~�+�e՛���	2�wG/������:�vĀ)�o��33؎*��V����������C�$A��B�<�h��*=|IJ��2�ޫ�w�����v���'��'G��׬6�-���Eh`W�.��Ü?�}�.E�|Ç�����>��B��&��9D&@�0}�Af��B�����|��1��! pg<J�֘�U6%e�+F�v�7���ݹ~	�i��4�AߍK{�c�ȭߩ�B��5�O�]���1a���k�-w a����_���W@`'��Y�~�}���?�u�C�q>ǆ�(��L�J�
,��O9�D�2��>l�D�:?'>}8�\гlP�3辸f��=�h����|����Pe�IM'�o��Tx�l��𡏨R�S�L���ݵn�M;N�M��?�o:�tyX<�� �+�ܝޏ��:Ďe�f��lw�T�6��4J��BA�fW�w���3{�Ȋ�U�J�I�|s�����ߴ$����g̷�ns�x4ӑ������b9�)�^�Z°|���"�|�eb��F^)�Y�d4r=���9�	����p7y�`s>��SͲ:KK��������x��!�
�g�3@w��v+���v��8��*>�s��X)�w�^Ivo�a}�Y��-9��I����+���P���-��OjB��BA}ѻ%���X�+�\��HA����O�B�%Z�Z0n����ǴQ�xoȖ7�d����{j~��BIlYܝy�T��$`B������W�\�ӈ����:�u����M��H��F�u��~\�;�ԑ�;W�4+��U�xO/1�OrPuS3���S�wu������������)W�+1�P�_Gvp�Z�)���n�.n+Cq��S+��՗��4�!:�k:;wwս����'.�6ʌ��(Y��@�0��d�pH�58�����қ`�~�ڋ$ˌ��)������F]���XU9e��y����^܍���]����#Ԡ�QI(Sɰ��(C>��4�ԉ�4*�̬i�.�o�z��V�J^��IU��MG^��E��)����^��Ib���-X����������)�<�ľ��
z�:���
���ndҋ�W!ب��6����s�vGpʩ�l%�:�'0\��c����1�y�m�c3^>Q�g-+k�y����8�!x"��M��yeHW%Ӗ�v�L��o�xQ�a7���R�剬m;�e^,%�o~+�,)��ŭ�㔭��K��(�n��~�`�ʓ��eܤ�v�-��%[�O3�6Ӈ���L��Z�rV� Q�J��έ�q�54�����Hy���{y��CL�{Q���z!e�M�ޟ��Gq��ݣ�,��Q-�w�h^8vQ.��M������p���v;�.RivJ�]��o"2���8�6��f��z?��[s��NexK��X�V?ɒ�t�e��(����,ٽ�o���&�x���M	���p��85M�0��S	�I�Kx��+��;���() 4t�h��&l�������jp}9w�A沸�$g�ڹ95�Qq�N�W ����ʹ�����G�&*S��o��/7���6I�H��M�]o��
�AT��OLJ�6JF�3ұ�IN"�:8c5�����精t��TQ��9���*�Vɧ����E]�� PK   W��X�7}b  ]  /   images/c5f41113-5d7c-441f-ad39-f06af9a8b0db.png]��PNG

   IHDR   d   3   ai�   	pHYs  N�  N��"��   tEXtSoftware www.inkscape.org��<  �IDATx��\	��Wq����c�{gfgv��5۬/��)F���("�X�+R!"F�����#Aز�m6���]�w�;;;�s��3����w�����O���.�ݖ�7�]��zU��ޫ�^�]���>D��)wb�d�����p8J�M��x�Q��iH�xڇe�3̣��zI��V��ϝX&��\���U�9��:f��h�P���$X�pbf�!oV�+��
h������i&�j�fJ���Q��0��� �97:�bН%)���#F�w����<�%*�V'��z��fs��Qxg:f	��P
5�����i�Iöi���S�o0y�����)�C�����Q��7�{� 3���p��ӄQ�PG�!�U��;�a:�L��	̡�߻�s2�k�2�	�;�����8�eH�<J�Q�"ux�n�`DC&'��`�0\�`�5ޥ@z�, a_V�i�B�=����e����qd|l������E�{:ZW� ��E��{(Ң{��v!f�?Y�������)wsǌ#��q<?�B�%�*����М��B����ᖫV���qz�O�T���L	���&X��^ӖAS��'φ��u5���˵�^�:nqî$��������ݽ	��fI1�M}o��!�v�8�v ����XN�7���1�<�䲻����%0���ଯ���z�486v�3C3��SC!5��jΡ�)�Gτ�1)o���
�}��Q���Od�b�Nʏo`�)�ߦ�eXm�ؘ�.��ߝ$'��F�%�􌏤t=�����6�`��[	�$t"f@��D�If�ҷ���Й��I������^"WXc,!X%�6M#��(��"b�;+�$ac~�c[rK�J���.��?�u�|h38�X��k�R�f���1ˮ�W�c��^Ni&�X.�*نd�K�,AzYU�λK�D�E�
�'=�$uWI/�F�%�ؕ�`)��� ;Bm���:�t������7#}s���D���Ӥ�]�0���ۚ9ƶ��y��ʙbO�g1a��!�b��o�E��I.K+(�ؠ�P�pV"m�M�M�QOjP��2+o��l�4%@ӯ@_�`3�-�dn�k߇���Ͱj���c��H��drVJr4& �t���	�'�u;������Qlܽd���\T�E��P�D#�9�&"��^�	�6U=a��(ڝ��r�Rdx��!���(�</F4j�%�l�g���G��w��[xn��"�V�n�S���,X��1��V�4p���t�&Bv��P�,a��*	n3� �A�4�{�}���y�m�h�#�����(��wt�&Lj,����,����&��6"�/���4�B�p�:[���#3����Cس�C�?ta
��*Zښ���$��S���mGMM~�h`t|K�q�j/�~�&摜]$�;��gjk��,�p��d����#u����1��Z�;��X+}��� �UD��W��u#��`�ܸ_}C#:;��Leqfp��\�����	~�|���R�>�g%���㖲<�2C4|�8�
�Ģ�R%���l��M�%�]�o��d��	��H��Ko�V�5d`]N���ʩ���P���ġ���IֺX,PZ��2Lw�|����@*�&"9*�P���JR����&L����U�A��ԖN�x�j��`�}�v)U��_P�.]G.WRmҏ9T'���ߔ>G��K�_�Z��TFn�p�o�M��ot|Κ� �t*'F������
�h�Q��ф՚��XM��K�Ee�w��9�7=�$�`0�g���<�BmiV��Ό
���C��C�E ��@3��Bx�0>9O�Ε��Y���qJgrg!�2����2S�o�����ĩ��*��R�X���s?���VI�%$��a���vQ�]�Q�l��W~���tn�qc�[����L$�B���-x�bi���� �����N��l ;щELN/m��%1dc*)���'M-��1��b��084����;�N�q��I�����M��>���<�+�&Hsش��%uLل-�V+GL������XZZ�]w���_����'�p:���[m����xu���ɞ�������Z%�����u��O�63���"�m��������ӆ3���'n;�mm�HҶ�c��<r����|5�UV�|m�k�:9!�M/�gf�h�D[��ر��BKf���dd��%���<v6���r��Ѿ��ؠ�B~L�,���w|�3x��1ڳu��u�p���ٶ��,f
;����Rf��[*����,�y��7�=�N݃sS<��������*�F��jIL_�������S�s�\d���=�C��`�LY��>İ�&sCG�_�닸��G������|wC|��{��lY#������S��u̷��3��1C�]�Cf���&Ƹ���?��]�+9��7<C*��$�.�F2M�By��e��/��LF}��9����s�o?�.4ԇ�9��lr�Y?�啛��ێ��%�%Mՙ._U�,�6�ȯg��c�V|ʕSY�T�������(�JkOkR�07V��夻��V�; Q|�t۠�������(��ne�uy�:K~$�����o�:i	g1�⛿�AW�Mi<p��*a��.F�.�ZBg
z��x�/#\X������W/�POL���tgwCڒ���̹_uy�J3�
.�dc����ئU
۔]�)a'.[�����zJ�y��Sg�w�eqxw�4�//���L�d�t�^S�&u���C�꼁w����l�S�P�:����V���|܃唛�*�Huu��S_bWJ�oL��*��ģ���>�V�8�>O�������n��c��ӆ��9!�}��/h��c�rN��li�E׎f?y�޴�ӋXX\�C,���	��I������D"]�������*��thW� a5ľ�;n^�(#��K87�ώ��:� �O3����������o��_�^o�� �M ��������|��9O�L��_�w|���G߇��>bPZ��q�¤����j2#g���`����� O<����0�����<�����u�a2�����MfO�[ɠ��Z���S�g�3r�~����ŗ.���dp䅳��Ղw�z-j�|ph�iF}�� IG{[�̚���i�v2Y�ֆ09� G��\ՅPЏ=�;��{�M7�G��f^A�sYe�g�o�$����h�S7Y����5!>�|�]b+�6̱Cp�������VM��A�0��3���~�� >����} m��8sn���b��S������8���)L.�֫,���R*�Q��b�:1Ad)N�B�ňo؇G�|ѕU\����)Qao��]�z4�u�"���BLȡ���lC1켨���%��.3g��<Bjk�;���݊���T�V]���ZA�/���Gv�3��n��:ë�'|�$:k�djR�=�����f_�x��uV�RM��5�J;l+N�ˌ��3��y�lۈ���Ɍ`f2sy�����I�5��f����u�)�3���o�&vܵw6�=�p�/z�qg��n�^�sn;��XKj���;*�)֗S�e������Z��՗�Nx�{t�5����U�I�����:�d�{�� �E1�LM��e	6_�s_�.���W�L�h���λ������M*]'՜�����ǃ��O�^��
3!�+��<Fj�g�f�`��p�>��>���y��� ���7ϋ�2���5��͠���o	�xjU�d�����u��� �mwh��O�����+���]�;���j�q�����a"�W�Q�R��g���|a�[l�����L}n!Vv�t���k�z$���i�V$2.��mf��VY��Xd�*_T�\m^�jȞ@�&�~&�����m��28;p�--�����S����h)�yѠ���r�U��y+Icf��qo����=Q�U!�Wބ�ZKl�x���ބ��(b�8��owbp` �@ ���Sr�w���jo%��K5��J���ϊ��nI�
�3rE�kz�c]^��$/��Ey/��y11>�CC��|H�i	~��W���Č�]��юK��_cؐwv��ҒB�z%��.�PЇ��y���������;�W�]C����7�n��KM���'�����;W�0艧^Bm����rs��sϡ��7�r���En.^n��b�K�tPn���U�Ea���M��~�-�ު��iټ����M^�b	�������x\�`Ng+��pb�1�NDԫ�-�e<؁�#���'`��m�\N
��3rH�ʤv�k��H����񤱶��v��&5`Xul�z��Y�`��꟫���G�	&/������tխSG�o����m���6e����>�ۉ��4���G�mү�򂊗Y�)�B��+'Fpwo���W�i<w������߅��Z���3Y�85,������\�wp�.q�O�,b|rA}�v�s��%��oO'��=�L���:����?o��}t�h��؜<.�r�!�n/�i��>,���xF^4��r�Į��]��������s�s��ӄ���j���*F��RG��/Z	���=ޗF�u�^d�"��3gǅ��a|��ߧ�[��b�)�Q���(���y���~^eXXYB��Iĭ�|�`���I:�f��+�����D���-={�/,��cZ2�$lq9A,R{%�J*O3o��f��Nb�I��/�^���ȬH3�V�g
>�OpD���.��0F�%-m��T���r<��Ub�z�-�+���g��$p,�[̀{M�E�2�8'��-l3d�	����)�!7R�]�ɁD|	�ļ ����`bb���sI�K�4�#q!�a�h��[o��))ǁ���U���e5妁�H�F(�L@sx�r["6�Ċ������C,�����KF>���*�y���ޟk�o���22Ɉ�a�R��,]�*r!YD<�}����1��>L�1h,��g��D�dB�1ᮤ� �?GDP�+E��H����Vy���R���6n�yЛE{m\�ۨ�.ڿ$J	��9�連)��@$F] %Ag�eeM"�p���`w��8� �)�j���ql���0v�.��l܏�d������.�f��9ڄ��hJ`;ڄو��&8��S4T���`Rpb��,�֗�ߓ�%I``cZ+�E*M�m��J1ֳ�2�8��͕��fH�̢�;�Z�#����q�1b�	qdP�:�!W�Ys�S��80�S6��r�KĔ�Vua.+$�n�@H����J�S�7�'PD�`�DtuH��ƣ>�R�C��� �0��5��T.�х�!�R�M���c1�<u�nn=�Q(2���fB��pq8𘄧AL��Q|�.��7$<��R��M��� a��z�����k�۩�����o�|����l�WgZ�眛�єV����2¤�-�7KOc�.Y�rT9&�N��s�F�2��2��)<p�N��%?�1$��'�T�	�Wc&�N⡗k�-ZoΉ�o#�/�D@�0�����^��-3��p�R�f8�U�9�{_{�F��)���а�9+���p���b`+���ٰ�&�1��ud��S�"�<�0G,�MJt"���@~��^b����jl��J%C>C�����,TȠN�����D��χ�s(��[+�i�d�T���OPqY0V;cKLF��rr�鱁�2�$��	_y���-��,��c*���\PS����G��̡��0�ϯ΅����Ϗ��ݹ�h@چ�G<��S6��YqK@a�5�(1��ӢT��d���OBE`�G���Ǳ!�ɏ,6r���]f��$�ӎ���3D7s�2���G\k%�(G\sav���}������k�f�6����0�;Ov))1�x@���۰:�J���a�r�yC!϶��b�hk �dG���Nd֢ޑ�X*���^�.kE�c��ޱ�d|�g�D�c)ZQ�8��4{,�������L�����a#8�}�t�?��q�d�    IEND�B`�PK   ��XK숤u  �x  /   images/ed2519dc-d5d3-4f03-8887-20886b87e6c8.jpg��eP@%:8,0������:�n��[p� ����;�-�m����j�ի��n��u�G�����Tu�-�m��HHK ��� ��m�� ���/�u$T$$DD�w((Ȩ�00�ߡ�cb�����BGO��>>>6!.>¿�HhHHhx��x����	�A�#�3F�����!������ pHp�5 �W����2
*�;�� x8xD����_��_������M��7C*<v��Tj��.|��#� �w�D�$�hh?��sprq��򉊉KHJI˨���k|��26153���rrvqu��{�
	�O����������_PXT\RZS[�ohlj����������_X\Z������?�sxtyu�������� �����?>����(�����$"�G6d\�o(����Q�D�r��Ш�(_�9N�# ql}�������P����F��y[` ��[0��E%7�3���p<����%�B���[a.����@:�)��t4y�\u��r�ƅ�i��<�f������\�����C����	��������/6v|��i�����%gΪ�<����]彩Ց���������Nr�P(�~O��1I~vs��jԵ �8J�_�B�y!س��_���[u��#F6$4�!���e0�� �4iN�6�\�ۢ��fTT@���T�L�fw��C�,;'�����S?������wd���;d�b�l�klI��*O�
�d���7 X��
���|�A��CM�}���G�H�k�|�&��^�N�~�}e��[�_��t�K��"�	��0N���Ss�x1>�#f6�}jd 0����r�𔏼�p�c(5�k��NJ �rh�Q���8����,�x���J������O(�����F���C�Z��Oc�s��em����R'��p�C.`��i}�ZG�����'�L�e��� �{��M�bmb���nU�����B>$������Xc|w'�W�)�:�2��[z)�D��|�ZS����Q-���o���U�������:��zri�iٟڍL�Prex�y�c�t*�Ҝ�Y��	{���6>��������͋m�2c��ja(���7q�yJl�m��� ����?�F�d-�������Vʹ)��qjqGq�|��Kr\Q!���T~:����ˤG<���{�%���/�^[�$P*lQ�p�炘c6��"\�C�Q� �m�P�	L1�cp�i�>>0�\�˿��0�K	�2�1A�~���ܞ�\=sVI��!w!�슬����-Ȩ72��@��j]�m�&�x!gu�|��cb�kJ�|��0B\��fZs��K��	�IB�o\�J�5�*f�H�E�}�{�w7t�lS5		��R�����޴����d�/����A� Dv�D?��A,�����U�ٚ���ś%E��`����N�åŔ~��AD�+�V��˼i��G(u͒�f�ӡ�f0�UCts�6��h:_K�y�\�^�+q�E��/x����#c���)ψ��������]l#�q�ʡ�����~C�u������W����Z���j�8B�/�MR��q����V�
]���!���%+�����)m��¨��j3|ʽUx3�X8��C}l ��R$��6�����{%6�Nb�Aa}A���Os�C���`B-V ϫ T;�p�w�s?`��=ݙ�Y��>ю�w�x���\l�Q��-�h2d��m�[�2^A��y�G�6�qz�I[>(`��d���e���� �Q�PFTɠ�p�Y��28�19Ӭ�F�a�(�}wR'�iv�@(�P?<���.����B��a�d��4E��/2�:@rP-��h�:�G��#2M�L�r[�[�ٮa0[�-�8ҹ*��g����]�����s��|8 Qb�L/��<pH�;j��j�-�4��/�YlyY ۴FZˁK����H���J^$;#:�k�m��%`�z�N�B��_�?v��c
A8.����T'��;`��T@O�zL
՟���J1-�k��·U�Qw��i������Pe�3B)�J�����d�;!H�3�"7�7DVIi�K�-�j
�� �8j)��5���^*�)v���s�=��x܊OɴB�
<�w~��6�ڴi�(��� u�b�7q ���E5�*���_���D�F>v��.Gݴ��
��N��tG^�R#�)�K��¿8?E{Q���l�-7#m�D��T4g ��̎��c�fۇ���3w�[��į�N=E�Lp[]In6��3Aێ�0R_g�T;r��a�{��<i�_�lBŖJ��	����s�G���&���C�2bZl�a�4�ԃr�E��%�n��oj��ncj�� ��/o������3�5A��1��}Ɗ���D�E��j�zE��� 
h����c���� �+���i�@�U��a�=�Gc�I���Da��;��Sހq�fW���	����m����({28����:D����Y(�ʢ�����l��K����o���T2��]�F@��=���9%P����,��G��8?bQV�>Ʌޱ*M�q�W��}����Zd�����p������\mj��&c_Zc�!-�p=o���]q\sSk����df<7sA��f����ŧ�e�氳e�<.ܭǬi�l��	Ŷ��(�i�EB~ȡ<��չ�A�:�ӫ�2mm��/�۽��H�h�fL�+��7�E>����  ��+��
S.�L���d�dF�q���O�l�Y��C䛿6�q���nϱ����+�g9�q�n�	Sm(A�޿�G���y��Zis 5�c[L��8/r>�u�Fv�8������q�����,�Bu� ءd�|��f�7v^���\镭����W&��~��(J3	k����Q��~�O .��e|)+�X�8��
y���S������@=����,{4+�i�X��ɤͶ`�S������*�&�f-/ŗ]t�6��\��O9k�I�6�(P�����{֩���
+�%��X�L�̜�֘����A�J����(�L�Gi��S�>�S��Bf�/+l9�ڻ��;���� �t�-Y&�*�Ǌ�����Ȉ�5�a���1�8��n	�ȚнL �6�7/U2Si�D��gL�S�����4�a��S�z��n�Ӷ�"��M����r��kJ����7��uf޼�oW8$/ߌeLo��o�|6^L����.���� ���M�Cr%Fo_Z�Ej�UT}��5�R;�^wX�]��ne��O3��@-�|��ޚ�h��9�8B�-����(�b�k��㘑�����M�I:C��Wj��9�^���ޝI)�u�ݯFƕ��:�ͦ��ҽ���#f�Y���f��O�b�͉B�L��v���,�{w[F�[K͖V�M�"Wt�ӕ�R���m�!['sk�7dl.�|&lږ���e�j�I"�g<K����C�|y�`OUŒ{��#�b�F�tawk����q�;�]0F-�A�c�ZtG�\v�~��/��m�-�3���5�g�d;ʗM~'�sƠfE�v���ߦ��|[v!���u��S#U�����Ȼ�v�Oٶ}C�;9l_�c�����~d��#K�Vb���^S�ć?$o	�Vm��,�ǳ�KVq휾�U�rHy�E�����˂#�E��%%T�)

̋Q�D�!���m��]zf���ͺ��sL3~�Jr'���ʟ^����ZYBBg�ʣ�PB�2~����Hxx%�ܿrN�8?C�1��rv�W�g��6J>�x��ߡ;��Kc�цԉ=$�g��2{���z��S{�57M�Y\ʗ�v�e��+��ԏ���g�J�ER&�T�_$	"\o�3ْ\���hz��\!s�c�)�0��@P����9󭴕c� �м��Ǩf�T*Q�/�ev������-��I����4���r	rR$ȟ\�`��eq������_{�Qh/�����WTb��FĊk���LM��mw�Eg$��SE�{в�t�]�P��H-Fs&[�i����͌�]����z��,F��sk�,��ɷHW{�pj������	��dǲJ��P\�j��<\��(��v&W�v�ļEy�i�H�
{��l:>��z.�a&�b$�i���س��RG֫:j^�м�:��׊4��5���oj`#{�ճ�ה��oG|�æ�������-�p=�
s#b�k�P���_�v.�?�g�o�%�H��/��|FW�H�� �;J[+�+������V��p��K���䣣��e*~��2���R��M��'�#����ȋC%PO���'l�}ٯ[
�o �������'.�_�\��g�Q`����gyR��>�K6 r��G�J�W  �	9,_�D�*y���9��� |�����
3�g` }���k�pw�����HS|w|9v��t~*A�Z����wh�xM�?�R�%ט�|��>|��$�f^�B�c��B�^b��%�r9�뢠Oיr	U����ͯ�T�(����+6�A%e���C��a����	ko�v��{�RX�&[�G��J�QG��񋼐�N꨺�h�_�;�b(8�V���4~��z���zC��j���O�]~U����Uz:�m+��H�X���S=�뉰qc����uU��/6�E*� �Y9�t�r�D`�/R���=��5k��v��;���$H��}E=��Ys�X+c�v��+��^[PM���J��%�vD�!��Չb(�Z�}/B,���[po�����9�
"��i.�Ӈ>B\_�%��1f����\�݌���H�O�s���"\'$9��I�:Ps5>�?.qΙFR�_���ى��,11cz 1_L��d�e;�$�-���9�1dDu��5.6���7�h��ȶ��"{���c��OG�F�>1��� ��4j!�h�dMj�ɨ:ϰ}ʆ*��u��?Rz5�!�������u4�/~�1s;�Z���=Q���޳A�N�Ā�+6�~w}_A�{�o5�|?��q��B�6|�|�?�/klƤ*�f��g��R��m��yA,�*&w��-����s��u��L��-�����:0�9�����\�꒗��ќ,8�:���y��!��p�d.����Qpu~c�9)���<%`���#�e��?wN��,��xTq���b_��RD�G���]�i�9yG�E!=���Zp#�fM�{����g�C�C[vhӉ.�v�n�F��<��k:�-쁍^�Ȋ^Fy���܌V䔳��@l�Cs�$��#�
��N\�n�G�N�Wb�dX3q+Ks!��D��/m� �eMfz_��5�(UG]���1���[to��`��'	�3�6w<~ c ]ldUlά92��3�6��a�@Om�������m��/Ⱦ�׊���jI�݋o�lye�p����`��$]�5��>�t�:D����N46�s�{c��W.�tҥ����5��������\��(m����O2�o�<�V G��K�=�l���'�%��"�����xyAS�H�� wn��_
^%l�p� �\f��/=�OSfSiIǴ�+y�������URJw����������;�D�q�iS�S�^K��m��x����8;ZU��v�zo���t���0��a�G��D�[��.d!��y޳<��,�n��$�Ք�j� 7�ڐ}{��
�Ⱦ�����ڴ�Z��F�g�t��	w��Q�Hx�ſ�k@�#��`@o�iu�&B�n�L� 5J�0JNy�͔<f�M�߻Ϲ��x��"WM����H�\����%�x��R@���~o����/��g\,���hf6����R|Đ�f8�.���E��b#���sμ�=ƶC�ԑ�c����8E��Գ�5/c�\EU�p��tCò�΀��׮%lc��}E����fV�=�9�(�{KX�{��0H�m7I?�-�8��L�s��j�j���{ �sX�S�8�e�k(��˞-��+q>����d�� 7�֯SW��qPsC�؜�>���.^��1��Ep��3)+���!A�u��gn2�BG@��}��g��������߭��g�D�߲
m�V��3�X}���ѻ�Y��=�����$�5@�����(E2�E{%��m	�.�u�D���_iC��� �g�ޜ��:�H�n};ǴyS������D�k6[���'Ix뤓���e�<K+�٢Yj��RI�F�J����O�\�}��#,����y0oъ%�Y6�MHl��@�ן�$�@E7k�X�kŨI�k<���ZR�����E]��ӿ+M���8wdޯ��V?+��bQ�p�ٽ0�0��Y��j,��� 
��~�5��p�Z� ,1�q����L��N�zm��c_3�Ě��a����y�*vz�K�X�	�;�Y�_i�Mq�%l#�+�q�x�?�g���6Qv��� �$�֗�O�hi��M��djCdFVӶ(�4v����枆!ޒR�"6��_$Rx_f"����jl�,UsdR�)k�����C����������JjIaڟ_c7�a!��MU���z�\�}��'�_A!�r)�RD1�����/n�ZC���0o��k�������/��(�8,�H6��A�!a�!����,��
%�g7�0��y�y��7�?7�2IZd/mk��kz�[&�4���g�ߝL ��"[X�8����������M��5��Ҁ�h� `'���Y��0IL���aܨ�ӓ����Q����'�L�&�L��g��m��ì�6���h�C@���F!_�<RCy:�]�Ȧ�J5���_S����4to��f���k��{�C�4��O�?W���"�P�p���Id35mab�����;��UE����ݭ �^�^y��Mb����>F�3�ïJ���9���-��5+�P~ %?�
����۫h����]}����̹W�a�ozP�9H[�7�9{ر�s�h~�=���yE�'e!.�C\��$��J������zXh<�Q�}I�Cj�:�݇�^���ޭ��y�@�w~���U�Kr�5AP��ܪ��2�x1����Q�쎮<(d$��k�St��I�����W!��!GR�_Dj �U��5L����/�w�lг��fĸ?���S�8�:�<��DV"L���U�@,,N;e%i�#Zr��`��������y�T�Lߥ�Bd� ا�ԭ����5�_|� �>�^!�\R��CK���:�����Xw����͓��;��Q��+~�1���]�+���U�2�2�[1X9G�q�J�%��%��!�l����³���ˋ�i3�ӈS�h>n���OW��l��rld��*J�E���f����n�9VJ���/ty�4�_A������1���U.�8�_ʧ�;4�@!F�H�VS�����Bc���J�&���F�0��y��QW��<S�	tg�_캫G�-�"I*��,ǒh��)��?��K�1�m+Zz����Z9�w��&A���v���}$��v���u�u��jI�����������tm)�;�Yu�˘��&�
#d�gCo�>�r�#�O�mb��\5i����Z'�����L*��W����;w�N�whCG-�r���$],T��^��ʇ\<}�����TW�m�7B�H?�WO&,+��B=�.�p۟����dg�L�>g�h�nq"� 4�ӳN��2V}1��;0�M�j��B��6����oL��lXiŷ|�'��t��lr=I [��1$%����q�W�KR�u�R1׫��iwҀ�v���TG�ǵf���%�Xz���ͪ·�":kZ�p֋�VK����JɻJG>dJ�J��K��3&�f%���;�$��?�"�.27�zB�R�.Mm7c�i*����>����M�� �U?X#q4�4�+��>:pه�u�9;�ƂQ�\����L����:5��VrV��(�����'�^E����q���i+Dz�Z{y5�ƩU�� �N[c�u6RD����}�H	tIAD���kkn �#$������7��{�7 \C��)b���$���e�Y�3Z������l'
a�CƊ�¦d�70�΄6��F����Շ6Ar�|sʲ������$�K�Cҡ�`�黜�uᚃ���1sn�`}���x�3�h�B<��r��)��ظPkA�b���|�3~���Oz@�T��8!�Y5�
푹������ ��M�R>1�D��Q9h���s[�>�P�]���YAx��m,+��G�7�^L��M���4�"�_�x2��Z��O鞤%������&}�^����?�k���.�
��_�_B�:��uT��V��[
�g�j-=t�k� �cO|�)�y(��b@�H��a���W�bh��}b90J���NE�QO����HYK#�i�x	-�^xF��":҄tfhY�rE~Q$�T�f?Y��7����\�����%Y�T-�Ū��՗���	�P�%������������J.��A[�è�}�t�qWq3z���Wأ�
̈��vH"��-��:�a7#��0;���2�`l���hZ8��z��T��ќK-�k��$Ϙ�)1�Q{�*��t���'����(U�!r�vW�=�#	3�IéE�j�ϲ�u�d$��fa���)/�Bi�[nU�m;Oܘ-�T��]��b����d�_���س��҆!�4Sr����g��GW��9L2��V����C��4���_�.�� ��k�+�ﻄ�+�*���j��য]@(��4XL��V���s{@�yi�G6�А��t�ԭ@��- ��}$� uRm��JV��	��)�*�`",��N���ˎY��Ҫ�����N�U!|F��� /�3"ME�^˃y�~M�j֩�Yf�Ɋ�f�-�2[WM����t�����;�8B��/ʃ�Ӛ,?��� =K�������aB`�o��A+�נ]��@�3v�y�\Z��@�o"غb����c
��+�F���h:�,��y��,W���J��=�6��R�vEe(8��@Sb�sӧgS��OĖoܯ*̾@�-�$��f��E]g�j�]�Բ�t՞-��q��ĉ;���p��E[�r{��M���oU �|���I����7@E�!�(<��۬��s����T�Y�Ʒz��W��%ĝ0ܯ����.�=�rY8��̅W�Z�W.�?Kփ)��\�b<�]3�ad�o=t�g�s �ga[c�߸^�G�������wê�ZDK:���VC`��{��縠���}����ؔ������4��pid���
Ia��Y����+�5a��2q��L��pN]��Leu���A�"lY�D$'	�I�����!�+��D\[�x��=���즂C�jY���~�Ǐumqj1�37���H^6?^��Y�g�������$�x��JԷT���������� ��,�t�,|��g��޻��j[�h���:~�R: '�����}@Ŀ�,�f���n�R��b�m�%���" �	�6��L�I.�j	�����a�
pD���%��|�#�N*�/E��C�hu�Q\W=ݏ6�L�2����1
���Z�'�rW�dk�]&�G;�8�������S��l����9�j1;4���(�{Wo�]���U̖��F�Y��q>d�~J HDD�[Kg̛�`���u]���ȏ�L�ۄֆ#r\�����a���Qb7S��g�h������`�&�VS�t�A�e/'D��z���
g���8t�.O�,9�t �XFA�c���*�˖��x���|jo*J����6�'��u�e/aFފ�����L?m�x��6�.~XYT[�[K�&�Hqs����9�6�ģ���WX�ȟp	p����%NC�U,]љ��e�T� ����,#cd�{���x��������ڲ�[���=�˫y��2l̂�h�q��z�>���z1��R�2W|+�m�Ȑ�j����B4RB%8�}��ԥY8e]9"'kd�W��kZE�뿬�s�}OY�:��m<����2r�ƞ�b%̒���B�.�f�Ȍ'�j��t�&��:<��_Ż�p�}z���N��ɵ�9����@`�'IJ��l��x��B�w'6�G�V���#��%���`p?#\��<����K�`�t��z���Q�ӱʆ�����}z`�e`��]��d� y�9hL]��w�<���d�E��$���Mۏ��suc�W߽���	����-�UG�h�'������Uw/
�����xpz�^�+��b֜?��H�ۺg�UP� ��"[`6�0�sƴ���]�V�8���㮼�̊kj��Ԓ(x��՚õlƪ�ta���W�����%��j�Xy��C�$_����p'��*^j-��ɑn~�|�x.��i�'z�%��uU����1���b(���O�1�C�V���B� Y��,�NGIͳ�d�=_�z��3;��q]�#m��[���]���ͫ�o6�'�8�H��q��ծv��e{�d�����}���n2�j#�����d�>KjpR�"B�A��q��b@^�^Hu�\�,Ѓ��^�G٩ނ��^Ҳ�[�&A�Å]O��P�WD��)Lq��GR�1Z}Қ�3=!� ?u��6,_�C\]DS�{����E%��#��]8�?@�ڙ,�).^�=�TS��՗7�>��:���ţ	��Nfkl%�ו��7��~��5�NU���A�$u�b��pA�~9�� C�蘫�W����(ؿz��1vw��JW�����8� &Kn��Kv��dW䓶��k[x��$�.^*��6[�B^	�*�=����N#��d!��Q�?�?�_��_�qZjp�y��wn�U�ah�5���[he�y���Ƽv��^���I�/B�XEc�q+e� ���v�-H0+&3�jj�ƽ�QN2قy�V2N�Z���εP(VQo�[%Mj�y��EQ9���%����*�|q�l�<���i�\*Ih�8D��chk�{�� �=f�Qd�~a�䮛K�.�uJ\�;�Au&�	���p����(r+� rj�������������B�v(��x6�K�1wh3��7Ib�%�i�cgu0�~����]��RK2�I_2�#1�ODY�V����d�Ð}�����.�0!�xYm��)d{��t�E���OU����t���i�b���c�m,=FT��<�p2�]��؈���JiSe%sL9ڜz��5��W=
��q�����L��c��84��إL�2R7�����e,AU+V�+{��{�!<`#�q��}��J/�K�_����nM��F�JV$&^@���nA��%�>�r�"ӑ�B�a�3

�TW
���ߙd��,���Cd-��K�����s'�s����?B�S+
TR���B�F�Ǘ'Bz��Z�~��I�Ŝ�I���2�ɱ{�����S0�� �)�η�����1/�D�|�V���m(m�$�Je���*��v!��� �C
�S���E�L��uH�Wh#^	 B�6��7@l�t/�ֶNݣ[�Ia�Q�r��r�����^2��u8�Qq�<���Q,��gvE�w�4(����7��(K�ىە�8.ҵj�q!H��$?ze���9��]c�ctb��\�1����*��!��S(��R -)�R֫D�ω��8��A��v*)@-�g�XbG�EN����t~��^ܤ�A�Vp�8]�Քy{R���3�2,��o��^㛤�~UP%�-�:]�@v�*��~w��v��J2�8	����3^����E��=]Y��Y�_H��ࢤU�d��ԺL�n���;{9E�'�FX���`���b�W�8JF��,����Ґ��b�����*n�7
"//*�}7~z�E*��Y�2.O��v�c��	u�э��ڐYh�j�ke���ݱRX�B=b�Q9��K��ȿ��0X#+R�Vɡ]9ǘW����߄~�׬���k`ڒW�P#��ݪ`�������Y��U�m�gvo�����..��tC�=�Vy6:X������-6��d��D��.Kqٷv�$���I(�n/�sɨ������9�,ձ���ך�����gX��򷍡OP0��"-�H���.�DjK �HfīJ_p��ڀ���8��>c_t���&��%δ�Űi� ��!e3��50���5�����5u�Ne��n��	��C��#z��V����u������W��ϔ�)�����8�B[?��tC=��կ��%��?)+�c��G�f�;��Z�}\ĭ�6�.^�/�j�#��m��7�ޚ�M��`qU��(]�E�����R�5�瑋��k�؞��ɋ��_g��d�Ar�s��,b�=,�Mk���Pv�%��v1�Ĥ�%�a�AU/�f�V�8S�z�O���s��Y����8x�缭����DsqV81��_c�����M)AD��"m>���y�t��9�K/3�R4_�L+�܃k-�D����vY���I5�t)O������ڲ��R���i
 ��E�F�������i��Jf���bܭ�I������e
���q�݄W}o��-|I�Z7R0üH���I���ϟ SuD��Di`�4��l[�%�$��n��zg��.$�J ����p3n#0S�sv}\��\]��4��\��A�'m_�X%�.����@��,�cs��@m�vg��aQC�r�4\���+1t�Jm��D5̃\<�S&ﳧҷ���ƀ�$�nG���/�9��^������I[u*i��EaMR)Aҁ�y�jx������^�����~��a�����k�-�?G�Æ9��n�q��)�>��/P8���zI��.].��W�Z0ݠ����ֱ�a�Frs`U�9B��ȫA��I*�p_K��c6��{�(����c������&8�}��T�������M��Mⲩ��f��7*�\V�V�bYZ��~C�r�۳�9\�D�럅O_�㄁=� ��ga��#�b�(Z���Y`c��[�1D��Gu���i�@�ƎiJ���1Ϙ���{[��E�wo�8T�Z�<�����.�B�J�5c�Կo�H�eR����|9��.��h<D�_���6Z����궬�:�fG��B��D�aܭ��0�sk=�i}���&�1��aJ��+vc˥I���K��Wg��!'��� #,��p%!�g��\/�����(�Y&�E�L?���途�W�Ɗ��<�H���6��Хm���a L)��*�0;�%䯞��ﹷ�H���?H����MP�%��$��� Q:Pԙ���hQ_*W�O���ۮ�6�U��3�r��ݏ]�l������ܷI���D��E��+p�'.|����MU���7��ھ���Xy;V�h�s��}`����հ�^a8�N�d��l�G���A���y�" �q ��I#-�w���p�p2������T�jG��%粙t~�Y�j̡S�K�W��7@M�Ɂ�f�F��\���&e��@b��e4֗:_l���"��F��CYq����u�<%F�O\���e�ۈ�����:`P�~���+Bm ��E�x�	wt����Xf^�%�"9�ֵ�>�6�t�7̳x����"$lj�#�b���=�f=Lg�zo�����%=��,�?r����@vz��$�T(ђ9��HZ���l�$r�O�ItǶ�XWO��i>յ/Y�5»�C�_�A�a��s�G��xF��S� ��㕮��\4l�M�[b�ׂ#�`����76�'�@�v�]�+V�u���s������U�PZ{&��z�2��W��3b#٦!�Ez�7��v�$�g&�z�+^�y�)�ңn�ʼ�>J�8]�B��:�ҳ˜�~��$1��hͲD�!�����UK��`��(9������T����rk��d{<"��#�࢏�p%�p�ԧ�5 ���x�xeB��	=�_~2�R���`����X4;id��Q�#��H�
y�6��|1i��_#��/
���\qt�ֽ�����#�U���Z�(�
]9����"5��פ�K|��!"�[�w�ըx�{�ɫ��hM�%ǎQ�n�-�T��V?s����"��'*|p@���8�AP���֋�&�	���G���I߼Q�fz��`z⻨��׈��k�dl�K��s|I�sǏ�������é��e���Z��鍭ŃG!2�{f�N�$�y����h o�
��\�Y�����٫9R	D����0�#9�
�aH��@�n֥��,NʹQaS�Ej�D�×GZ�p����H�w:��z���k�M�et5��}�!����F�ݜ�].dU'N�U�W��[tt3����`����SF�秪e����^�,�����M����$�O�*���+��6��S�T�����LK���9�{���+��2�z�[!4u�+��)ޑ¸�����&(�	��u�a<4>�e�Ϡm�ɔ�-=K�fu҃�Վ|�&���`�T/���O�W�:\q>{jZ�؉�nL�[�"���
�_�����µ�ړ/Ǔ|=����ڧ��L��W�	7��P�N9�DE�l�z�J��!���Gʠ�=h������)ةQZ��MUS�jv]�֕��}t�t��!1��71!f!ó�d%�n�4��I+�>DDDb���F� ���7���Y�º7B�}b{�k�l7e��\�%��x�}��o������K��%A�w���4�uR�ŷ�}4�H�:I�J����"���0��U�i[��B�Ȳ�
�~m�jn�M�1����̊�!G}���ˡv�{)�|	�K��%Q<�*���Bu�o
s����D7O�=�E_v�[�`��O�^z�j7~�_�h�x�J9�ѭ���Y��`WC��Z�lwպ��0����㐰��$jM�R��|��`:��{D&��@�w��A�,B@E����Օ�xM�3ƃ��k��5�p�(���?�v�9�нUěC9�ؙ��tb��M����>`�@v1�d��7=d���k-Te�������@�$ftZ��Ի$ǈ�$�{�q�p�6���>ס'�5̶���}�4$(��h���M�ݣຏ�Fo]#���"� �Z ʚ�w4!eC�n�Ny`m B���U ��p�9P^ƒ�g�M�tE��ٳ�9϶k�X��n�T��9��@��ܶ�����^�0�P��Q�M���|F>�Z���� %.Z��9��qa��{���;ٶ�7�DSll�v:��t4�N���k�j&�=#��½J��6��P��є�lIvb���:M���KE�K��/�(�؊҄y~������O=��G�����V?��<�7�� 3M�N���^�+ٮy�ݵ�� �Fq��nmL�Y�輽�p-1�+��<��WѶ�P�F�o�T��9���o�Ҕ��B؛ӰR�7�a98f=6�q{?-�����\�V�ZeLN���Id.gF�1*WJ��x%���3�^|�~���-�f��W!<�3��x�8i���h��>j������*��=��Ea�f�ι
�R�w�����/
������vJ�t:�Y�v����ۚ���4�F�|h��ģ���FJ!$�L��˾�Q�6i���F��j��S��Y��rvA��S2�G���όܥɔ�v��]z������o�tb 3+
��ǡ��;$�z�U���.�V��K]�$Jӻ�>�Z	���IQ�@��v��Y�+�X�{5j�t�S:�Y�ںQ,ٕ_���B4VA/)m"&�i[�rJa����d���� ����]���h����b�l1�ny?fq�J��޴_�]䴻/i���"�-�t ԖC�A$���{ErB�*.l�3/��d�sv�����B����z)=7��+�]�<�Ґӿ�^D�h�L���҆��p<�Y���o���O*����77B���8V�XGBY���X� ^�ퟟUk�E�Rl�� 4�R������OTH7��Zv�I-��/�֫�G�����?�$�A^ʞ��wJ�A�B؄Ba^���F#^�I��MB-����U�.;I*�*�"S7��Y�v����31c�&#�yB�����[h;��
��N�����\�h�F�����g��j���ȘsR�H�'�O�B�ޚ`�J���n.��Ϡ���,�~�*���N),-1��c��9��������~B�;?ӹiŗ������4q)���[�o#^r+|��C�pV��.]��jg�Sm(��?A�'?�B���e�������q�m^�xu��:e���k�C} 4��aMGO�b�]��Cƃq�CF-�믽��y��(s�F����;i�#̀hY�2�?���_�A��^�;����j����l	.B�
w)<��]www�[�����

�@�P�s���}q��t_̟����b�%�Q�eӞ;�'q��+�_B�Ē�Q�\>�0��o3��{����|���|�.`x�N^������S�V]����<��R��������	
�`dqe��<O�i �dOSVV���!v�
@A���)HZ�8��B?�T�zY
�$P%�m�)k
���ӂ��lx�	eT�M(r�g�n�5ﾯ��|���'��%C��y�Σ�`����ے�ړ����OB�j�]6^*+��d�a9�VU]h�`��-Nv-�e���C%��Z1�2 T���sQ�ٱ�z��k[� ��`��6x.r�V���<����3��.G��S��(�)	>O�.�������s���Wן�o��;��>}!)�I����F�r��A�HC|����&��G����`�|����w�J�̱�V����Ĺ3�X��&�x=�e�igÛ��#a<(�Y�����������H��=�C�\���8�����3KoC��N����(m��	��&_Ȳ�V6u^E=ۄH�dj�T�}��Q��1�+���,6�d�'�1�e����]����0����LiX�> i	Qv�Z	��%sbq�¾ɮW{Z��>qo$8ْ��f{)dA"'���ϽD}�3���7t��߯4����Qӯ�/�^�겋��D;��pf��2���SE�a�����bV�\��(DV߸\O���B'6Z)���-����u�P��_U�yeL�d���5I�q�#r<DQ�'��^�`�=���������@GB���:�$FC�T7���b�1W.�4F�)'Z�	����沧N�*T��Ó��7��py�L�ԭ(�����8��-8N�N��.�GU�瞿���M���>j�]6�������*��y�����Y={�˸S��_"T=֛��i�K����/@6&�>�v�!}��L/|퐬���Y�qq�H�4 �f=
�9.S�� �q�nH�ޔn�ԟn���=Ŏ�������-J[+_�v�A�����}�R~�'����|��gUnhn~H���i��MgF5S��vVK-HT��m�<i�ހ��۬�,e}.�:7��OM�H��MF��h󉨓����яٻG��/)���P�=�z8�%�V��*��MCFU��ed?-�5�k9��.e\��E��#ΰ��(߹N@(���E���o��[.�ڽ>̍��ց���Z{Y��:��s���5��r�EK���R�|9����}�A� ���BXe�m&Ξ�?N�б�U�ܸ�4�/�N�h���d���b1�xQ�c7*�6.6�̽�q�e� �^�z�PX��*a5�|�J@�:����W�g�h���R!ƻ�X�>>�U?��G?�K����[-�n'�J��1�`�m.���w�;�H����g0�֡��5��M]hsMZ �֔��ju���ah���������k�<+b�=�jq�� �X �k���<4�M�����-�pa�/+4�u)O����K��X�)9a�6� `�$+���~On��RI��N[Ɉ��"���+�gq3y��r%�S`+�����zD�E�a�y�Y�t���C�S� ̽}i�q���֤�Y��ϫU�3���fD-�*�Ga��Ɏ�����ڔ���Mm���y�
BZs�ȣiu:S������^X�E @Gh(S MUȏb���6��'��8B���3������O�Z�';%e�z�������.�V�)�o��>>��4����D����s�҂��b֞�}9�>�u#���ե\�������|�'_1U(���D�t1�n�]� ^�s�d)�����p'�L9�Ad�r��L�q���P���9�O���~y�P�c���b��?���M�j�.������i�m��D���[\o�2- �$�[��L����|�Z)�ӥ�r�qTh�f$d<s''�{�Pj�IqvwR�A�Ƞ��7v����2�@�ջB������c~��Ui&�j��6�͝�h��P�@*�U����E���T"�V�4�y���z�vư~��==�(����i���a$-��G{�on�Y������)�n��G<�0�6
` ��Q�۔տÿ�$��U.%/��e��e��fv�7.d�'����"W)3?=-%���A����Մ�<�Y�#4��,�ZlZ=�	��Ϡm]�z�]A�B������}�1�<Yg͜��"A�!�SE��2�����m�(��'.��G�Lމ��?�͍��KC^ɠ�'��07��%�]�G�F��<��|�{�L��TSu'�������`#�������1˾ZY�&8In0�r�V������^�O�+�`�!���|� c���岄b���撃2&\�6��xe�S�?)y.5�$ZS�-�E&�ǅ,"��#�0�}��X�v<	���뎰To��7Ga��j��[EX���"�2��'�[�S��A�����X�as#煮,f���v
x��Y��>�Y���\i]��J(�i���.<�,���M�śd����!/N�G�	&�F�D�]y����.�n=Y��� �����.n'��;�k�	6��]&#h���8���X^���/����i����g�>\;�v���,�����_��U�Ř��XpN}bHV������Cvq���m��YIra��9��.'*����[���Ӕٻ;�\�D�(�uޒ�N��?!���P6^{��ynOOc*���6��.�H�uPT�I�d�e	w�m��Br>�X4���ə��k:���b�!v�w8I��$�z�4���.3���j|-Y�2˞�l�_���T����Ae�a��y�/%�~�r��u�v��
�f+`Py�.$�B��a��8i6��<ZLf��hƋ�,[�oe�<����:��//���&`��ڿ�e�+���"�Gɇ�1?�����C�=�K�j"k�,vg'�.k	���q8sWN������I��1V��� ��W�	��W����Ws:��m�{Җ}�9[4�\��y����_[x��C�������ǳ��F^�b�JF�|��3%0^��	 >�j�gB��I�X����dr�^8ka�īxr��E��Z`�y��(�L�ٔUq��Z���Nf�LN���[��#wݐޢ��%�r� ��'����N��.�9�ݩP\��[߈i�q���5p�������%=6�G��W�P�Y��L������勇����:�ߘ���&ˤ�^3�H/��������~�@i�v�y���$n��_�����6ǎ��Nb&Q��m;r8:�5�<�����>"v�\���_t�tT]q/��E[匀��q��5-K�c�Y�c�ㅙnRi�4�y����Y�s�;	>N��}�"��j�Lk�紴�QRm�3�}�ݳ�@��D��{z�G�V���Z׺x]Yv#���3�?&�n�*�\y'������vn����l����D�Q�9͊O������4�2���q��\�٩�j�+Q��F@�Y��������iL��C�}��
�f}�*�5�'��?�=đ�F���������jW��������f����~�t�2��K�������4)�gE����r]��k.��BAwS$�nr�S��s �e�o����u�/��pq?�+G;�&wv�����d�֨F>l���P�VV�S�6�؞��Gx�>��Hxּ�^err�'���lq/�����Y������I�X���he�e|��	�o�|}Z���� %j�����G`����ix���;�J\;��x�+�x�t��-���-����51V�j=�/���g���xo�G��<�%���9�C%��z��do�<w���0��']	�&M=�g��I��3�T_��X�Mww�*�Q�4�x�/�)ֺ?i�?U�P�_#�=�~Jo��sH�ypM��?�7 ���TMd9�?�2�� ��T=YJ�Bg�5z\���3c�v��=�y��t@�.�ގ�q�K�#��-WP颃���lT���� L�*EQ]x_�}�X04>`׺tEVGWڂ���c�ze�ۤ`IߵM,�8����'���@H�����t*m�^��mɖ�1�t�X� B�n�8���i�j�U�O�����m�Aq����ISH6�H��R߶�����#��OA�9Z��Fl1���b�(�ek3䛂)�c~5U&Ѕ�����~�ȓ�Q����2>��
���EZ䲺;~�����LE��ا�[�Q�̕�@��m-���0^	sH���󢹀+Оyns�Xh21p�B��p��Q�l��h�k��Y���;l���9_��|<x�Z�0t��%3�����|���)4x���q���+#хCzS4���b0D�%��B)?q�ϊ8I.!k��3�����a�WRo_DD�44�J���~E��.^�_�a��c�.l�jT�r֪�F��go�}Xlq$��g-j�-?��l�L g� ��&�Q�>8�|d�*159�y�c*��`��5V�T�ޣp�џ
��]�QB��o���4K���P�J!���q���d��qu�E�wU��N�rw�gI6ޖ�j}U��vvl�~�'��}�J9�����s��C&{�K�H����C��;�١�!�������y}iL�\��6�ī��E�`�1	T��p�h��,g�K�5p�0(����f�њ�M�wh;������+a�
�f��-ĿN�'zr�Q��*X�ˬ�J"1�3r@���ސl���޾��r<�֋:͛�>*��z��@b��v����z"Hom�qW�?$�UGԺ$q�ȱO` B���IY�B��_g�̩��L�1�R��8B �Q�U<�	گXt��8��.�3�<��N���҂�9���IFg\�4�W$Ò���<�����������T�5M�_ʎ�e1Vi�<���o/��y�H��.G�b������]�{`0��k/>�KYM�g��n}�xЪ����"E�{����E'��i�g=��I_���cs�p� u��q�	���%�2?���#� ����ĳ�'.�� 7�b`ǳ������6C��H	�;#���1,��C�(�=(`�w����-�++e1i���%��o�Y?��}���}?_�6�WS�fO��s��#2=^A��J��Ј� e����V�{rI�7�<~���
�����5����]Sm ;�^E=9���;J�5�M�|J�� ��cY`�Ie�C������(0�[Q�wnU����i2r0�	����G"��"�d_���gx�\k˒�*�#c�n�/s�D��#�H���Й>�j��&0'40�����L�aq��=�ץ[�3����[�䅶�q�+j���M��}Np)B�2��c-c�\,�b�F�i.�����-��WH
 >�.,�gQƭ-�	��Qs�Q�GךA�u�f6��$��e��Bm��wC�_~M�\��&��&�Hr�֠>�6�=��޿�:x��N]�mS�z/ҡz&}�i�?�7옷-���4Ys֮m�.�em�1�ś�L$�(Q2>����'�l�00W���\���4�>��,�p�X�\WK�<��w��0����&�z�b0F;;Ӊ�;���(������<�dv���U0&XR��6��;vF	��.��#<[d>&�֕��
.�8���"���̣�︴�u#�>Jr�^NYq�ۆ�"�k�h�v��N����r����~I�h@{��l/���u�򈽁�R
��p��mD}1�+M
K���HRJ���T�H���ڱ�)0�u�݁N�y$t��c��q� 99<1�Mb��3�k�N��NA�Mg���=���G�����G�4%�í�e0K��p�dS��K�5�L����qm�>r�����<��N޲�]`;L'Yq��{���\x@^�vy������pټ�D.U� ��0FM��Q�� },-�˷H_N5#4�}e�I
��]��kKY��k�v�a��|2гD[�/�⧮f?.��F�+�6mت�l�q��G`��F������z4Z��ʊS�Ĉ^n�6�y�uY��Jo�|6A�]��N�����%/e�&�6�R�4�ֈS�8i[���?&$!�Cp�"�${%?#�5Z��?�� ʠ�U�=��&��[���ȇf1#�c��x�M�	��*8��|[ົd���1�<e����#��1��r� Nq��fLH"�ݞK�W?�m��q��bX'�DG��K���}q�J)�e�]�B���oӸu�`�0���Òiӓ`����gHc=�N:��D҈�Q���Uה��Ʉ������x�}�R�-YָU���Aj�C�����rd&$��2�G�o�s�t�;�|�D�a�kG�r���7��,���)��-4nku��<���4n��� K�`R�&�?��䱢���\���U�3�doLB������P��8B��u��$Dl�OS�j�QK�b�[��^��=a��.�]/,$c�!�?���q%�������b�U3���"�=s�
�ԛ�Č������Ѵ�ኸN����iNo��~A.�s�6�C�l�Q���}����\�^g�b�6�=��D�4��U�j�j�vi���\��>��N�����O �+�</�F�?�Dz�}R`7�(.U���R�[���7�����us�eY�9�>��U0A�ϡXP�6�CW=/�8%��@��oqS��_\�|F�k��o��:~{��_0�Z��{����J� ��� �&��'Li/�������F�D�٪�U�,:w���Đ��B��X+�t�lE�=Z�\�=Ь����r�#`B�N7Ӷ����`m�3|�F�V�KB��k°|�� 1�>l�sTl��ڜNm�Ǵ`σ��A�[A����ƙ��Y.���7�����ܰg�l�"�V10×��T��^��+vϷ�o�3'�A�=��I�k�����ք3v�U
n����C�;1QX�0�.����\�H�?�W��$�n�U0�4�˸�:_S��1�5�f���%M��5ճ�x�$�z0��^�H^�7\T�uq�ӻG�5WX{��Nb���6�F�pʗ����A\1\8weO�k ߗDp�%�|`����S.���]݊��:�5�;����X�(����|u#�;�'�%�����G7�$
_2��,�2���l� �R��N���+�c�b���D��sj�5JI5P��k�$�n}�SJ�~��> ~�	
	R��K)Y�^�'wFьN��=�x��O�DD}�����Ig�v'F���q'��W���W�2E9j��-�>h��b�˩�;�葵����1��,�q��}#�.��A.G��.�"�1���^5t�G�a�r.�LE䫨�c��ecz_1� �òe:��}��a������C����$Q��N�b-ϑA��©�q���X�WN�;�cJ���!<:j�°�SNl�t�/�d�p#���;Ș��:"�~w�}��_������AG7��E#^j��82��e��`�h����I���t�*�"��`���P$������߬��a��W�{K?���"�QN3ul �?,3�s�Z�e0�'�������~+1�; �`3�H �n ������мU+����v�V�/��fX����EQ�^4�
��ƅ����T��K�^al}ϛv`:��5�yL�I(v�їt,v������l��8����/�Y^q������j�,�9��vڍÆ����C#'l��gk���/߮�� \�(P<�鋕V�A���~�7�<C��ʛ/rV�`i�ﻠF�c�j���xy|>m�J����e�g����ve�&��G<h�:f�}
�(����y�ׯ����'��4����:\C.6]˨T-Hw��y��-��K��	8�/��g�F�i�q=���.���+B1vn?�w�B�8&I^4�͔�S�c!s^*�`ӓ�5����tSx[Dm}B{uc�춾�P�P�^�Dy������wŮ���%�ӣ'A��φ�:}ϡ�1w�C���*�v�6��9�<#!e*�V*q�7>&r���6�
���qks#֒w�K�
ķC�`�g�O��|_7��Ļ[=��e��y7b�?�=��q�"$L�ߵ��`-0v��q�yARH+�*���ծ4Kső�;䕎1j;��p��7<LQ����(�5FW��*�޹.eb��RXk
@uXp8;�9�7%A^�����1|�;��E����3�s䢄�AЏ�>B��Vq�����]��q^��{���`C�y�\(?��k��j�аz4�(Ҥd� Ƶ��l%C�k�GY��]��H��&"J.��p{�pot^�@{�<�r=�n�a������jV����Ɋt�v�����!�[7�
�iH�;fc ����YV��Q�)����J�������?�iG��6cD�����7�����I:��㋸��X<��w��.P���+/[�Dz�qn=�j�X@�y�	u�LR�r���\��ڮbƯ�K�	�q�Xhw �IV@n�^�I�P��>]�nAi��I���a�t8Q"���SR�1 ��R�̤kaf��~�G.������IFhΰ�K���{��V&EW�%'�&ۼ�K�E(��[��!����G��N�M^<���.�⦵����.��+�7��&�kA�?���4�*�!�v/���i�$���K��v ��Z~|Z���荕�u�e�WU5�B��Qux�5?��+���%��@�VY�VP߱�-�e�ʆ�xR�ȗY�F����+�u$��N!�g�Ⴆj}�����}��5a���<rDyx�����~�k�l> ߴp����\(��Q1��� 0?����}�h���Ω���I6X3Eu_����#Q%�M+�<����\HED�Z?�`r��Y�eJ�2��?�3�Y}hp�߅��D��*X���>>���-XY
�CF�q�X�&l8�|�+i��Q��D��'�/Ŝ+ n��<��C�-��M� u����K�59�2�#��맦����)SF��	�g&�Wt}�I9sj�uV>�Q%[�9�V�3���$T�J��s�^�CXD���%�ڜ_�X7�q�<�N�Ѩ�	�q�]���z�btD]�YJ�zƟ��lna%Uف�� l��)���i]�'�}O�D������`M�lҶ'Q��:A:9���(A��A-�#���!�s{��7�e�����=F��Tؕ#T��u$�6�A�4^�,�=���n89F7�J�N�W�lے����wM���!*��>}����d�&I%z<_��e	N����	..� i���άuG�:!� ���M�tkQ�UjwdK�}��짦��P��F8������~bD"V��\	y����ݳe�Y> R~��A}6�Kr��7�㦗�Wr�s��~:��z�k9���g�;L'���=����a �x)��F$^-��.^�M�p�AP��r Н.����|�=ֳ��e�g-ym�
�ݼ�nK�jO!;��W����?:���ܶO��d��Om7zn�+G3�*k=C��n���y�o��h���{1��v�O�9#���Ô{������-�,hl�ڤ̉��t������M^��ֲrW�Vb�� ��~C*�䤤�qڶ�b|�]��_��%�Vh�Q����5��He,�}"ͤ�v���p%a{����ǣ���-�)J�jSb�*��f���I�z'�	�~w�n�h���b���n���H8���IH�{��R�E�t�ϾJ2U�f1���P��^��i��8� �dR�c�ɇ��z;o����-ǃZU�Cĩ#Dvy��X	��5I�,�/YL������ ˤQ	b\����e���n�%��f~}�\���=΁�S�4�$+�$����Nwz�����#4��o�����!q*�w�Q�B՞܍�1cN�u��־>;F�� p1�[��Ɗ�㳨�Ԅ�K�>�,�@����Z�yEu�~ڥ#� ,��5#���g�;�d�]�Z��"kn�]��`�M�W���SL��������&�)*/683��AG��q�����2�����4uXP����dM��a�O�1�d�4䡕��`���A�`�c����<���w�u��@��W&����/�(
�?��1���'�dQ�,���Y7e�܂ٸ����B�6W�*��6p��L�)v�y�ң�|����2"���g�\춽y��ܛ�N)�7�{):��i�nϣ*���h�K+T�,����~E��B�qA@L�:_Z�Tޛ8NbJj�}���>j�/�P��`m�i�&}q�(3�mc�<p��!s�F�s�+3�m�����\]f=9:�"��$�Ml�;�]�b��>��o4e���J����tZ�i6P�"�`���H��Zʹ��5�a/�U���W���3�bL�@��4�d}oJɋ��?&��M�õ�C����t��'x~��, ��r'v�Ab�'������1��^!m�ow�4e����Oa�JK,���I��-��	��1�>�ں΅�J��%&#�Y�}�0V1`����(��DV�Р����� 	;��!�FO~���S���~��֍y�X,��&�+#Dt�I_����g����s�Iĝ��(*�"��B��ٲ��|ù�}�2̟ ۠�sKX1t@�����џR�az(�8
�O���sS�`��ߜ�{0k�6D��5�ev�i��[6̎��RX�tڍI�pmͪ�C�Kbb�Ə@gv9�IA��m�����"F�~mw���֏�=mW'���>Z
L|���I� ���o��b�
^r�6}m��3����C!�ӡ�<�Դ���>H9G$/T��JDJ-�뚣�a�_�0�d� ����7 �u޻�����u��"c|��R�R�~���S��دh��_׃4�
�l���l>&@�;���H}�<�R _��-r�2M��3����8-�@���F����܋�la�u
���y��7��j�t����*5���*�����?_��է'���;�bW�a�2^�^�i��C뙢�"�n'�έPOq4.�c|��<AB8A�K`�; *��ty�s[����ٹ����\ ��3�ܨ`��Q��3t�C��F�I{�.�������Nh4��������g�W���F���]r�Ps�����]�EPl������d?t����yv����[~�J���s�Y�Y�����ʱ�D� �X�-/j�|���I�T��{�v����<~\r�s b;K�N� ���a#�)re�>��Dlghx��i�V�`\����m�<*��x5��$;��)���7Kx����h�]	��ᑥ��l,i�Ȕ�@��e��gӎ�d�<�0Z���iM
�TP�Eg���Fa q��:�62�4��v	��RA<��4��.N&ަ�����|��-1�P��Ix��>��V��K�Pƛn����}�H�/N�'{���鍭&#Xݡ��F���7�u8��vC��8�mWW��I[�P�ݩ|�0(���`ӭ�sjD��E�����X�������]-��=}o ��H�ݻ]Î1��a�����{�=����yȎ���n��{q5 2�ep!���"�f�Ч/�ҙDR3C��=�E����W�.Ŷ����䘒�ˣ�e�j�Ͽd�G���tc}�G$��5�����_�L_���,(A##�����	�a�:W�GC��}�^�;���pi�d���>��hLp�*�&�1�2���{��g��f{���,ݔ��K*�:5��V�"&���	���{�����+<=q����t�R����r��";ͺ����A}���Є�3g�|��X_6�arQ�|%��-Ϥ?��L^H�ȐcA��=l��9����sCF���R N��,�WՉ)Cy�A%��=��}��(��#��&�]{���y� W��o�(
��	�=�ޚ��h�?���xƾR�캏����� n��^X��i��T�����G�g�I	��O�9I���~�AU1����� ���qo���P.�s�X����A�M�� "�Г�����@��Ղ��=�f�5���c�+<I��� Pz���G��&t���&�]�����kaw�m�:/w�̀M 9HM�^[K$��;'�5Յ�o&|�k�Y���=M��P��O�#��;�mըl�b�
c�6ȟ�3e'�eSfo�X���}�p{��-c�%%����'������$�!�<{�Cۏ�ٔSv��mIx� � �g�u�KN�4�r���-�Y{#��Z�ᑨ�+C�F^��u�!s8�Q����q< E.H�cK��n#��uY�#�߹�G���"���O��
I�MV�����X�a��x�1��|�kC��6�w�͚��+	e��P�D���]}(4��3��o���k�'��n{��N5ÃK�$'-�ݗ�a���D�Y�ԑ������y�jH4XWm*X�����=��@��s�M�C��`�Ue�`�i�mI�Tu]��CDAk�KA���1�,�K���ސ���RQO3�臎aңg6��zڛJ�r�cF�ş�5q	y`�?ߐ!�:�4#�鱝������P��q�G�z��Ɨ9!	?(3����Q����sH9a��9��y����)yEs^�%+T�\��*�9ѯj�n���)��:�̯��v7��!	��[0	X�;p����FK�m���Me��֕y�
n�c#��]�r` 1�W�+�|�R�,2���G_���ƫ6���N��jJ��F ��W���`�q���%�V��pɓ*4&��n���'$�Wb>hi�=Pm�P1�T6��;��g��G�8L���{�w��..&�PvV��_�Z���ކ�Sp��Y�>d�0�o� ����,�P���A7o��H��u��~	 8��o���T����gA��/�Z��?���҃�8�%����� �~{0�_%�|�Ƚ#�\��<�Oo5w�C~��(d6���G�� ,P�߳71ŴI���7����7u��� v��YNߥDс����QXB��Y���z�H���I [��m[>u +UL�e�]��c>��i��X!S7�Ym�T�uo�<��~
�Ђ�aJ��<�s3�t��Բ,Z�{��iF��j��Ěi�y9蚻x=,��Eu��W{Z�$�G�F�g�����aNB�����`Ѷ��=N2���%�( �U��Fj���>|��<���F�'��|��@=�O�*�b��N�=PD�~���}��%o�vK� ��-~ĩ�S���qR�Y�m���l�-���:�Z-�����%���N��.'��n�?��4%��Q���7��'��Z[������+��T!�8�!�DN��{g�[�or�\S��5Ikk|q[�Ƚp�&U�ޯB�wz%(��cUྭ�?PK   MP�Xm��c2  w     jsons/user_defined.json��_o�6ſ��3^��$��%�l�&AAQT���<�Y���$�N�'G�~�.Ϲ���rw��ˣ��6���XVu,��忱�VMM_��g@W�wyw�vy�ח���m��y����8��t_�xݴ�t��#A'Ыղ*�n# �#�:����9tLBp͵*1����G��.�����m���{���*��^�����%'�U,�`����e
L��暞�T�i]6ˣ/������n����Y�;.%ϤF.鶧�>4���ʤ�R��"wu��m�>-�wmU_w��nh�U��w՚���6C�(VB:Ȭ5��T�7u�iZz��e�>��#˯�i:����G:�������W�[\2�\�T�t�m6��U��wG�z(p,�WV�B2Ur�,���sk"�P���n�:ֻ�G9�n�u��!�����O���ؿ뤶n|{�M�k��:�)B+�+�/��K�P*fs!YpZ9�<H�s�|���P��X�������,W%�(!���f��+�SE]���j��QG�����X�<��T��О������0%hr�� �pA[)3��#=�ʌ��~���[�@4+�e����E5��Ř.�&�DE[�C��t9att�A�@t�)+�}-]��cFZ�0_�T����*c��+�c��6�\j�EG �뿺4f�$����e����)=pܛ@\.~��]l�?�Vu�����L��j��Yh��"8f(��Aa�+�3,��F,[�R[
��]�!�3\D��K����>�3�B���P�b_|����;2s�����*��k��П�/�'�V�N�kP���!#��E��H��]R������Κ"�;��������@|��Ӛ�W�ݢ)7T��>��PJФ��J���4QJ�8��y��R�\��ќ�\�T���R� D6b!�(�. H��RP2_H��.���9/��N9p��L�)G�l�w�z�d	+��
�3�H�?@�r�9����N�95��x��ˏ����J?��{"�.�93йN��9g��hc���Ĝ�ȓ���׀Wɚ<�}��x�"Y��$i3�����.ab4�M�KV�۳y��pڻ�%������S�iϥ���Ĉ�C��|�|�w���S����V��S݀��Ґz��+��+������ c��2�?��`�a�Q9X���c����߿1.���ck�a3�_������öÂ�pI]`o��M�7 L����Ox�G H���0tI	����_`�a}�8���_`lb��!+��%>�9����0�U��.�,0Ń�9��x�L'Ҹw�����ii���~�\}�PK
   MP�X��Gq	  kN                   cirkitFile.jsonPK
   W��X�Rr5�  5 /             �	  images/01f582cd-60d2-4b90-a97d-c02e30bcefa9.pngPK
   8��X�bZ�b �f /              �  images/32499b6f-cadd-4b9b-b4f1-e31be966db26.pngPK
   W��X�@M��  2�  /             ' images/54862705-cc12-4a41-9ef2-e24c01e25159.pngPK
   W��X8�w���  ��  /             2� images/805fb750-7b5b-4a1e-90f5-2022d18e6d35.pngPK
   8��XF �.�m p /             ~g images/9fb635c6-6568-4694-b870-d787cbbccb08.pngPK
   ��X�,͓�u  sx  /             i� images/a2b075d1-9af0-4984-bc8d-fa1df8fcc417.jpgPK
   W��X�7}b  ]  /             QK images/c5f41113-5d7c-441f-ad39-f06af9a8b0db.pngPK
   ��XK숤u  �x  /              d images/ed2519dc-d5d3-4f03-8887-20886b87e6c8.jpgPK
   MP�Xm��c2  w               �� jsons/user_defined.jsonPK    
 
 j  X�   