PK   ��X�zG��  �K    cirkitFile.json�_o�H�ſ�B�*���~��]�f;��>$�@ITG;���N���SEˎ�*Z��4� ݎ���:u���a���d_��lg�ݾ����o׻��Z���C�_~���4�Nn���a7�u_�|�\v�G�?n�h��x��6��̔Y�j2�VI���:.�zYQR��*��yǳxr���tpw�u7�{����{��^)�F[vʺeቲ�DYz��=Q�(�O��'��3��3���������������������Lw�ey�,IIUK�.�<���*�2-��"_d����~�<�7�r�����2Ɋ|WQ�\��USDU��Q^JQ7�x!Y9k�?�����b�+n�����;�Ϳ�}j�Ѿ^oz#�nv�z�>�a;ߒp����!��t~/G�Eةvj����Z	+��ҋFz���m������Pi��ƿѹ�V[z�-=�Y�]��B�G���oT/�+a�OX�����',?�)�|�SV���O�OX~����'<c��X�����',?�+�|�sV���O�OX~������'�`�+X�����',�{�8tgQ�u)�,"ɤ��8�h��o��l����$5ʛJ{pV�����I�\+����|���	�X�*V?-?a�	�/�e�M;^[^j�S�b��׀Y��+ڽ�R�����_Gu�;:\ ���=� l��ύO����&��.��T}�`���R<>�W���`'J`+��1@4،b)vo�u؏ؐRS���{h�:�J	lK�)
LQ`���Lf��6���(0��~���L�Lj�S�b`W߀Y��&��&5E�)
L1��r���p2��dt��Nw�؞ �U������lW�)
LQ`��]ʺ]AJ��MO��'�c�R�b`���Y�m'�Nj�S�b`���Y�}#�Fj�S�bୋ��F����(0���/f����_u}�N��_��:�uRS����o�)�)E�M+�V�{vD�M+�b�U���V6���(g(^��B�kl:^��u��W�{�����T�r�,$*�Uc^Ѽ�W�I�r���tnoR�_��ս�z���/Q����u]�Y\iT̛y��"*������t^ɲi/p�ս�{����{uo�i����n��+cD&?��IpT}�D ��$J��dJ��J��TL�A��T�0�+L�
S��T�0%,LS��T�a��@�`��Sņ�b�T�a��0Ul�*6g��o0�E�8����T2�a�:E9�>yGmo�B��rHB���!H��"���>hG��H�8*�t��M�끣�J���Y���(=��A}��
*��s=pTP�U�>�G��H�	 8*�t�B^���JC���T��^K ���JC��TT��vX5���JC���T�ñ�'�ਠ�i?nG��0��$8*�4D�&�QI�3ɼ(�4O ށ�ԛ��F��F2�8�l$�l����f���,��yQ�ސQ�6�aI��+��@z�c�u=w�LxXR��{�������Qx�K �1����aI�1mށ�Ho�H�AxXRo�K�w ��Ӽ���s�F��N���L5/e��%��|�QxBV �1k��#�aI�1wmށ8h�
�y�#<,�e��F��^����5/���%����QxBZ ���Y��H�a��(��,��ض4/���%����Qx�[ ���i^�	K��k����@zc�����Òzc��(�q0�ޘ��e��ޘ�6
�@��7�y))<,�7母�;�]b��q�5/���F�ȃ����5/:��%����Qx�cB��Ȅ��\����}�] ����Ƽ (g�$�������0 ��y�s{��6f����&<�ށ0z��$J��dJ��J��TL�A��T�0�+L�
S��T�0%,LS��T�a��@�`��Sņ�b�T�a��0Ul�*6g��w ��l��	��	 �04��@Z(ҁ@#ݹ�ahTPi�t �F��89 �04*�4D:C��Jw,A�@T"��QA�;V�@ �
*��Ш��y �F��HahTP�{- �F��HahTP��a �F��HahTP����QA�!ҁ@T��TahTPi�t �F%��$�QpX�<�|�Qx�a�9�l$�l$��s�F����˺k�08,�7晍�;���f~0
K�9g���0zc���Òzc��(�C�0�ޘ���తޘ�6
�P �7f���(8,�7楍�;���i~0
K�9j���0zc����Òzc��(�C�0�ޘ���తޘ�6
�P �_���`�ܲ��k���0zc����Òzc��(�C�0��܆��v���%�ۓ6Ҧ�q�����D K��k���0zc����Òzc��(�C�0�ޘ���తޘ�6
�P �7���(8,�7母�;���k~0
K��k���0zc����Òzc��(�C�0�ޘ���తޘ�6
�P L v@ ���[��a^D��G9˨w ����a�(g�w ���|�ڿ�~�-v��~�^�>�.��O�}s;��ԋf9[og����O�߾��[�ڽE�Ïntg�XupQ>��:x��v���yw���|�L��I5ъoPJ`�V�į-����S����͞��2tz|k�j������߿�)���N?��N?�
��1|���~��^`�������q �@Db)�����>_gij2�}����P���w���\���z��{��]��I���F�?Q�O��3e�\ٿP�/��+m��P[��-A�֠h�P�U(�2m��E[�F[�F}.�V��V��V��V��V��V��V�y�{g��'p�����T��T���-�4%$�hFHSU1䨪�@v*���z�NU��2�ց�T5pz˕`QYƁ[( ��CDUS�rx����H;���٦���|�L9<DE5�@n)������ )����b ���CT�n$�RQQM1�7��!*��z.Չ�m_V���[V���@�(����9,@�(��������� 0~��L�q	�,C��  �%�������Y��>A@Fˀ�(��m?�R+���
%{����əgD��VZ����!�  #m�K�)��!?�R+-�	�,CI�Zi[�O�-gfJ��j	�C~%�h	�C0�P¦VK�"��%A@FK�%�Y��3�Z�m�Pb&�h	�C0�P2�VK��S!A@FK�"�Y�R/�[ ��O|�]�Bʽ$0�P��VZ�3��A@FZ�3�Y��+�Z��fB��Zi�B�g��Tj�6��  �%`�,C�Z-�mB~�"�h	�B0�P��VK��A@FK��Y��#�Z����2Z��*�6�`ҡR�hH��0�`��H����D�g,~�VZ�3�_�"2A@FZ�3�A@FK�3�Y����p|i�0G�p��i�w�c�pz'9j����j��Ǝ��s5�_��;�Q�������k����8X�[������ۉ۵�^!t�'W߮�ܥș.��υ�T�M�е�T\[q�ŵ�\\{q��0��i�]�z�ø��0�G��bO(��{�8�|жS�_�S�"�ǅi�P'��*uw/ж98}f������\�n���v�b@@���̿~�̝����2��H:��f��EI1  �_Vk

	�m]�M_OH����Ɲ���俚ÿ�R�O�G�d�����Q��?J����G��Q~�(wW�z��=���v��mַ7߽&'qo�}gO^Eu�Ͳ�*���Ig�fup�~��<����>�� �����n��aݸ��%n���z��L\^%���<;�15��2Yn�QXdW<?.�앋Ub���jUEI�ښZ�$J���Wu�;!G�K��m%Ӊ]m����ךc:������d���u���b�9�M��ʦFҫ�ٴ���Mbs则�6��LY��2s����]a����.���8�j��#Sŏlg
{�2.��ˎvb�vU~ԫ��k�N�T/�+[<����'yK�ʱ]��.�ǫʎ	������%����A��vqK�<�?�:J�V�UR����|jk�*3�Gyv�נ�4���m`䡸��C($���"��g� y�H��A��#�ⴁq�dɣ
'�!�:k����cH��!��Ǻh��X���,wpE��i��ae��*z�]Ҏ.-��>ifZ��dY@�'�lmXy|�p	�oO0�X~>�-׻�3�D����^9ΞU��W�.����Y|�Z�������lZ��"��<*��e�Je�ڶ��&�ҦL�y{�t�l��f��lzw�K�ܞ��I���ˇ�qq��~nRw�)���ĖO��ʘ�L�����U��2[FE��
�8��2I����N\]���^7}=&')�4d���4~�����C�g��f�8޶��a���j���?��ݧ��o���}���I����x�]�E��������O��ȓ�U��m쇷�����z�i�o��n�o��j����ޭ���n�Bǻ���ױ�|S���w[`('%�N��I���	%M��q9�Bꤘ�K_��<�Vu�E&M�h9��ԙɛ�W�����Q!�U�ā���G�=�eG>�X?q�$�t�}� ��ꈪ����r�ي��5��ʹ]�/s�tO�e-�ܬL3��b٫�z�D}j�ꮽ���2�PZ��~�u�n�vw�e[�ݍ� VW�����x{s=�Ū`/��%,܏�mOj�������]f����3�������ٞ��C����=؛}s8��˺��?�bp7b��M��������{�����d��Ve�?�Yo\��,���.p��w-Ծ�����E�w�����7������n�=��Z���޽�����Vo�?������o��n���̒<�z�.v��Vilծi.me;'��y7�b��y��V��d��qʐJ1cU�K�K�B1C
�-��f�S٦�VvU,'sq�4ܨx~�~�����s��+9��.9Tr��(��O]>o��F������_���<�xłm���I+��~���N�{�Z9=[�yK'�s�N�/P:U�ҩ�N���,���u���s�����`������p�VY,��{��7;ĳ���і�.~�-�AKg��G	<o�K�<�hջPF�O�+�{�?�#=W.ñM9�xڇ�g�紕�(m[efH���*�/��t���b�U�k�Ҿ�8l����e�J�]c�E6�Ub�7cəV��\��f���o��ٯ�ۍlk��f����o�����e���C����~���f���fq�ks�دo�F���?PK   ��X��.P9  4  /   images/3f03cad7-594e-4892-9bc7-779b63c9e608.png4��PNG

   IHDR   d   p   ���   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��]yp՝��{Nif$�dɲ����b��`s81f	,!v+�l�RY�J6�����M��&�R/��
7�@��p�����`[6�a�i4WO��^�屘�4�����z�4W�����z����!�x�	4;�_$��D%=����v�ho���#_��]w	i�8��C�y�h���9F-���=�r攐D"a���5��T�4�)�w��0'P�1V�a`|�H�񬣐f�0AH�!��\w�u��曱p��dr�n���[o!�����,�5[�*���:�����_��9�e4�h�MA�v��m�����5|>_������b:I��ѣ�<�`%R;�1��ӧ�54t;��6!g4INML��z�v׮]��	��f���^4!N��+H2]���n�Z���P ���9䩩��q��	��h7��{�p�P�GD�f�o/&p���1�6��B2m+&�mpL�I��N*B�Z$�jL W�ؒ��0�������E�*&�kl�9�$ep�&�����	�8�9��-����h��{��P[[�I�&AUU��� �*D"����6� �kE��FO��l�p8ظq#���/���B�=���	��駟bǎ8x��K9�Ԕ��>'�z�W��~�r�-X�h��8t]G,fFO`D�)�n���ؾ};^x���RSv���v��4�����R�&�>�%��4��_=z{{���9��amϗ��%,Y�dX2h+I/h	@-�[�:_�n��8�s�5�`������J�:[Bx��/�X^�N �#?y�$����EKKK?��{�x���P(�cǎqL����D����̶�|����V���生oK��ɓQUU��I�����_FGG�Y���\�W\q����~�//����������aٲe���+�إ�7ɚ7o^����9�� #���v�{�2z���Ǻu����E�&J�?������;)$�����w8 ǁ���,'h-^�u��o}�[���7M[ ���-!T͡�����ï~�+466b������ ��+M�E����N��;�uuu2J��XD�Q9	����/�555x��Ǳk׮�^�	y�=���n��ٳ��wZ	g�i�q�UWa�ڵRP6�h*���~X
ǎ��d���瞓dp��o�4}G*Ф��w�y���~7�&��A-x��W��Z�f��`2�}�݀�#�1/^<�L����-�M�֭[%AV(� �t�~��t����	�8|���<O�:�����r��̙##*���"���w�^iS���G�J?�`��Z�h��1�{�쑄$#+��o��M��V\\,���CA;��1N�7}#�W^ys��������'��~Fb9�!�Ԏ1ԩ��2��b��~�?�������<+B�9�р��*>3�s�7��h�dԄp gΜ��`�5�B�B�,s-N�LL.�^ky�BV4��L�>],�{:`�y���<��f�AG>���X�"-"GMYe�w��W㮻�J�p)���R�+ق��K�3w�I4̇�����[�l��{:a��M�$���u;���Q�x�x����N�M��.���%��ȱ7��t���+����k���jT�Q���J\��!Z�צfϚ5���7q����j2�^�Z&��Z����8��^z�tV\6�jg*p9���Y�dad�x��t��c�-RG�'��$C9�z��B�}*��x[�(�գA�&4#�/P��2�\�G��2��)��dP�R1Y�$���\�y����o߾��wF$���|uu�|m�d(r`ļ:��G�3'���8t��9�����aZ-E�Ԅ�Sh�O(�ӹ0,�E��Ձ�a��.8�5A���Yc_��R[��H�b-�s�ҁ��4SԌL"ʌ7�)3snb�,YO?ÙA!3�j|���at^FTh��	X�S�,�� P�?� ����c�}�K�Ku1�FM��߃ҏ=���#���~R��M�����֊Ć3�#����
�֠�Bl�FR��d�ӏӫB���$� {7|F�E�w��Y�����J�V"�}*}�w�W�ß�@�}�ZF�{E(��c~~>�:��$"+Y�}�\�p��x����^���v�"����@��?^�� �-މ�z#��N��$�4E�Wq�D�F��
G)ʜ%�;t�k]�jn�:C~f�4��˂�&��-!ӌ�E�s�!� MT��(�6��K"�fP�Č���!1p(r{c�oBP��ɳ1ɫ'=�V�(>�i��B�j�Կ %�|?_�-&@�2���(>�Jۄey%�d�L��ic�'!�Єg�������b�?�;ѽ�NpW�|^�SF�1�Є�[hT�����v|��)V�,��|8d �EL��{P�?��9'� 5D�1=��_�A�	���tĺ�R��8�.1�#��9'҅2�O5��D�%�xY|����pi�Ӥ�	�{��$H�)Hi��MS�B}F_�0S-2� ���x�����b�2"b8��:�����b�{j)q)�Uۡ��Օ�O
JCMŊu�3t�2>	5����I����9�j8����S/��1��^�B�(���K����ۡ��(-�/18�g�1A���`l�kE�5���:�R�@��V�/�F���|�=S�)!�CΌ:�X�4S�1&cP�R^h�+��jʅO����]��Qv�(��� 4��)��qz%�yMg&���7������4_/����U��2��Q��_����p;B�#�X����vh���!������{:$'��p��9��%�Yl.`v,�G��>�-�]C�v�utϏ$}�o�D��?��1��2��� s���a����~�dl��=+�X����9������,����l(k@BL$�L�+?(Κ��]Ctё���!�u�<�`�XAi��t��V!��I-��e��Ƥ>S�	�._�"�H���NsŜ�O�vX���Q�U��r!��G�b����"��D��&&w�h��}:!3�B'���#X�թAW�E�\YI�J�!<z��ؠvtǂh�v�jq0_`|:܎��ZP7�Nj	��%��[�%D��mWn6��{
N�:N��!w�c���c������5��0�=W�Λ�pBqY]/2w�ۣ]b�(`:$����S�t�H��-���hA-��o�M�"f�Px�u��na��8n��~�4v���F�A�}q9d�f���C�u�:¡+7(�'�-�B���[G� �ry�����r�9wꉤ=�.q>&x�J�ў�,�y�B��G�Ag��/o�@o�+!2*�D���㦈�f�O�P�T�zv_2�H� �-!� Qd�.7�y�g�1.�2��B��	2Va04ٗl(x�4DDUZX̬���ǐa��K����h��9��r>� ��'�9%��;D'!�.�u���ԅ��KP�ݭb2�4���кUٗlБG������t��~/�>���3��2�[8j�Ry'�&�b�8����0��f'�g��n?<M*�'��
�Uto�Ј.!��"�e�>X��9~^�i*��D�b����� ���Eт����;�wM|u%r��ə�[��L�w��S���(�@���h�!8s�{�����!	�;{��]��ˑ����0&�!�8�F���r/�K��D�Ƹx�b��Na�j�����t���:_�p���Q7ڗ��ׯ�r�L�ބ��b~�`�����s�=��%U(ֽ���m�C16�%p�4����tCH.����1�_I�eK�_)B*^s��)��GC��:��uK���m@R1��>���j�IE�^W�Ў���@�)�	n8Q�7��f�X<�K*Q�w�-!��$V�[��M���8MoGճ
�	D*y���qW?���dp��sQ���~uL��0����X�7���w����������v�ǿޏ8��b���Q��n~k+��Kf`�Qߡ�|��(��wB�骷}B#�Q��Y8���{O��1/N|M�Rb���P3H���<�6i�SUT���5K1���Bֱ_J��#�`5����A,��e���נ�`ڃ^4m�|%�>�>�۬��IAF�*o�Q\*�|uf}P�+�_�!�Qw�5���-
.�y%���m��tL���_��k��&�6a�ZԤ�����G�]3�N�d�2,k��)5��,
������P����k�e��z�`5��w0���W'�:'�H�`���P���������lX�����ӕ����{9�0��]��]�c�L������݈�DP"�����й"�pUB�Y�#�+&l$�D0�-��#�}.>ȣ`E�*4`9�Mʘ�a���i�xk�ԧ|�6̆��"�{`7zu_���J�8��#8/��t�R�G��/�05jf�E�5�.şZ���$��T�$�.i�� h�U3,d���D&��mB�"LI|��Q����ۇ8���Bqh1��b`i�=��D�⧁x1K4���Τ�O��K��C?UI	j��:U��鳰v�jTFʠr2Y�ʹ�9�[�ꡳ|,/��,l���V���+���j�D՜u8r�|�{?N�k�.�QŵX�-�.w��vS�&�$ȓ]�kԖN��b��,�G<�}r�a��d#)�G�M͓�b���Qo�����β��I�|QCC�,W���2��	�wa�g���SqbF3��G���3o:��T�3wq$Uװ*��	��9�Q�łʹ�+��6�R�in6�N@���q���z�VAe��袋2.KE�M�����O>)5#$���㲶�%�\�k��6eQ��/b:|�D$v̉�Z=�OC��>���Bsg+�;��`�*��D�b��7�.�]>Tx�Q�F��
>w����\��y��d/{��?�<(`c>�2�,��k�"%�����O��#\.���ƙ��ϞU�eyne�#����g�bj��+r�\���>�y~]~�=���ڸ	C�$��Ku©9���\%�b5�l��Զm�d�2V�怳�:K���~衇d�e��lg���ݻwK2XA����N�*;Ο�����<�Ԕs����-͐>x��vYE�7�2c���3�U#�>㩧��}a�\]D�́��(ɄX`��M�&�����J�ӁQ;�;�"	4��t�j��kv�d���q9��M��!;w�u�y2+�ߜ��MU*���5�:dEC�b��}��$�N�3�:B�e`�*8�H�fda��V�������Ê��`���@_z��y�M�+[S�@����[FS,
�h��ӧ�]�������q��!9�<����%Ág����L;��C�,0��icltr��p�#0"�������[�<މmʔ)���!��Y#��O*0�	L���2(3eO���`7fvH��8O��|�Т������[���;T#�V�������P��t�R�ǣ*(3e����~/��Z�HFV��dB�=�l�tO++Pf��>0�J+�Y:��.�����4X^|4`�Ĝe<�b�ʻN�8!K����29����TGY��o��f��w��Y�p�م<X�K�q|�$M�p뭷ʃ%�_f�7�t���o2�3�`Kנ��Яd�����O���{�DO
h]���W���_�^f����?z�}���!�\8�j/���9�J���S٬��C���;Y��%����9��e�:���΋S����ǹ�Ŭ��Q����t�T`_��6ȓ�g0㱁4��jE� ���8s���>��ma�ü�s�I�u��u�dr���V!~<5�f��1d���4a\�KN��bXB�h�}�v�p��*h�#���ߣ�;ǎ���;�>��;D������A�����5�|��̣�p}�ёr�� �p�ݫ^{�5�f�%t�AE?1��رB�\���{G����2Y��iK
׫�1e�N2<d]��{�����$��b�9�8_v������P�~/LR���?�G������$e&�K�D}�va������}�@.p7L'�9�������&�o�{r����EcM����邔.������%��/�ӎ56����݊���1�Ν����V&�Y�Q�^�����D�h���~�~0܋F����@�L(7\z������/))��C?�o��x�5�@��;�yY���>/B�l��+��?p �����kV���5t:�۝�0䓐��&TO��p�n�+۷ow�p�����9�%��<��c81��������f̘a�T4�+���r;���v&p6&)0�? �y�Og'    IEND�B`�PK   ��X�"{Q�? �f /   images/4321cb83-9d65-4877-9350-be2835182319.png�uXT�6:((����"� %9`"%�
�����e %� ��4� (�]
"HH���]�Y3���?����^�3{ﵞ�����Z{�o)�!;M��`��ݐR�`�uc0�?����.���Z]��}���χ�ohXa0�e�?����q��)kiuk��ck����0vvv�OM����?�6�4ǋ��`�1rRWo�GL�h�Y���Y�0e�@{�Dڂd�nA]�WO���>
���?��^��m��;��y�X���LK��}������q挑��6�\D���!�!�ѡ�u�G�"f�1�?�{�0�y��Ms^9���W���r�ؚq��hø�/�1m��+����`�LW�\��3��]����ޙ �7��]8^tv�B�3����A<�T�Qf'Ky��stgΒ�a$n�q$�������+�����u��0��_-�������o��{K�M,�}3L��4��������tU~+r��z�A�U�ޥ�����=�!���UֳQ^^i)��+�'(i�+�qG?^:����@_o([��}.F�+�>�n��:�Mمc���#]�c�ދ�{�)���o�Ӯ&]�?G�XC��ܯ�Zi�.���:�:���K�b�%?�TY���4��)�^/�ð��y\��Ƴ凒�}�&�zKXj�8[n(w�-dc��+�w�8�#s:�dw�u:t�[~wΪ��<�ϝƏV��g�2�9B�����@�J�y�}0G�lc����с�C�*Eⷿ��ӊ����(�r�|.m%圵��<��0������#l��gʊr��%����%Z_�K��2�_;����_{�h�k�=ϝR�u/��!����%^돓Z�S�'��*���x7y q��'��0���0��ƴ����!ِ̂��a���np�˚O{��%�$��Dr���8��}�*����OT=Tǻ[v�?��v6w4�8��@3��[B��YGjE��{��̼�uKVr�"M3V�tş�D�o�s�� v�X�T�b��a�O7�=�g�N���X�Uҕ�]�\c˷Ôas��ƨ{�E����(]3���5W�5ԫ�uv��o�s.��4�W�w� >|�y�� ��q֛��\�IW�vNP���Ф�>���-�Ao����7x-*\���q%�����e8~CʼO��d�ҤV\��]�}�.vC�X��q�U��-�����>^jv�!]Q>O�ՙ�ywϴk�T���!ҕ�DO`��ƶ)�o���0�uZB\;���ض����̿J��"����}cL��L�8e�L����.��d7ѿ�}�WF=_~��9-q����X'�}vĥ0��_�����o��1m�����+�)���1����yF����Q��p�RP�Ƴ�7 �NfE�0��+9�ƴ������G�#ח�hLUB<O������y<�7|�[/|�K�}k����K�u�G4���Io�eVt�7�S��1m��MzT������$$�:e�oRqEk�W�M���`�V~�epm�q�}L=��G;|�*~l�lǞ9��K%���õ��휎^��1�%��e��<����Uhߩ���=����A��&̲�U�k�v���}�t�?��_�k�����Z��f�#��q�ϟ?ͭ�Ԋ���	����;�KKK*ZZ���7��?~����� ��ۮ=��995QX'��4�����|#��L�lӞӚ9�~�ᗫ�f�m�/e4E�q���9��2��\\\��ļ�2��}a� Fll�)d�۶�^F���^�Fm��t;3eX��V/vv����_�)�9u�0,mccC�:`1�FVF^^~q�OG���R���4-����­完'ͱ���O��(��=�7Q�G��;��Xl�����b�k�ojjj�7���i�*_ښr�B}�Wz�x2;�'4��eW���eDFL�N�?�(.��(c��р�H��(�����SNp�?�^�|�p��Q���rk;��~�%�SS��at2~}����ȿ����7���ğ��Y�V�>ů��Y�uv�ů�G|�%)Yz�UױE��2�ע\�2�7�S�i:뽨�a�ڿ���a�|;k�{��O���E%ɭ��O�䱄�'�b�= ����ẵ�jŮ���#�^����9ɫ+aQ}
y:1�Х(����X��\h�dZmR�z��|l.��it�����,!�(6S8���`B�P�y�B�Z�%ZrOmk{J����l$K4JlL	����(�{�f�������A_##�	�W��<
������p5w��|(�:�q-�sV��_ORv[�}��J���(��C��N�}��=z(N>�;e�P��۾h�Hn�+��U�=�}j�t����p^��4�y�W�^�ZJت!������z�#����Q��Ήb\�"N^�x1%	�[��>'�� �a;��w���y� O����o��
�%EX���c�c("���=M�!��k�(�r�O!�/��pW�l�+�(-�FB��.����J����5��1���Q���@�H�#[���	l�A����m��H���)��J����P%���p߶󑊦f�#�����-���?��b1c�%ht*|�HZ�x|��2��F�=�6�m�T����dbb�2���г\{����?j:=�6��}ht�J�A1�����k��j�}� �444u����h��Q��MȚb�۪��^:��E�	��v	ٕz�ժJ[�Ĵ4�ⵟf�)IQ(y�����P@@uu�{`Ǆ��rm���e��R/�)��v3���Q񜟙�#�*��-���r�Y x )�ڶ�?ŕ"�n������#�:��8B�K�.T3���hV�ev5i�m$aUe�G��)�f��؞c����2"'EH��������*( �ҕO��Z�㋾�Te+��z!-"Ux��7�tno+IKKG��zS��;P��e�>�#���D|v�ed�7[�{b���S�8p��SPCgVH	@�tN��Mf��(T �Uh����ޯ����R&���^�;	����33�d������3�{����t��c�,N��w��a���g���;��@�u\��L/�p\�G����xR�ɭ"��GT�>����8s�t��ũN�╢�Ӟݜ�]�ĥ���ء~�rGg����iO~�R�SO��WBW�����/{���8�ȃc4�T剹=�u{Dg��qq�ђ������)^�������O~��H��O{{�e}Q���7� '�m;��U�&��b��Sµו����]o���̅�V�ϗ���Y�9�J�����3�wW����:���($��9��Tz�c�)�0t
�ײ�M�}���$�-�7��l��Fkr-�T�]<��b�R��c��?�����)X:L�&y4�O�v�h	U�35��Z�4�O|r!x��mMM���BD���1vCQ��͛���@hF:���zC&�i;<Z��Z�F���C��"��51���mU�oXp�0�o幽��㣮R�u1f}���hL��� o����P=��̇�i���iE�	� 8}����o�O����a���ڃ�S�c}%n�`j <�J��{��c�+�m��T�2�x�H��_�W�xd���&N�3�I�ik�V+�G�d�i��7��A����<��E3�����-��~��\S?� ��I�3^۩���{�;����|	S��ܡ�����<LP{>� |
¼K�����u�+�c>��~U|��/�}�Ŝ�Dt#�*K��Jo�;w�9�߸a�s��>�NK?�3��_X��� ��׼�Txm8过�7W��
�����P�jن���G�(ִZ�*�����f���%�F��=�^lJ
��a���� Y�-�X�وaH���X�kJ�*38����Eɢ��ecH��$��V��"�;�oW����4{��xup�*���\s�����O�@U3{�kW"o�R/����? ���mE؝��v"%I'Ć� ^z�p�QK �7b 7���B�G��!���/r�X�o��YR?}�YHW�
@@QB��n��
��J���'�wK���S)l��ϝޜ��G��;hFHH�XW��ĩM���Z�v���\�G��Qv��h���%$�>s��i�Й`�t��r��-)�`u`~~���X�x��r�v�{��NP�� 0��� b��z�/�������ye�B�YY��Bdr��ˤqZo*%�3K��R����6�mU��� /&]���䍻�/"�q�_^^�ȳ2�����]��e��餯�+HDp�
UPL�z�8�|s���Ξ=�[����h�u�]4K����ԃ�#����7��2���-k�PRB��D�� ��9��e��j����z���NN��t��������`�H�AAA�t�"@���  BxtBy�<T��L�N��ʀp��^�L��'�N�����9 q!!��-�o�0��9ȉ��f}��ɍ4��Կ����T�u����N9�독���`8��L���a �.�a��3���>��L��r��ȥ](��1�$�N�8����}�-�vG��׽�c��� �֗��6VX���?Y�rb 2ۧ4ۤk��?H��{����HKI99m�p6��n)f��\�dQI���W�CÛ߃-�A8�6��ph흷�"�_�:ޮ��Ǿ8���ｐ�62���{Ԝw?���]��������e	x�̹p����!��>���Ҿ�s�Us�3������<y��˨��Ql�K���j�<ٗ^#���V���Ac�$�:���Ko�w����{~%�>W�5y�KPP�W�6𤄳=��^"A��999!#	�F�͕K#��R|aJzz �*�4Hq!j��sg=}�&6��!�>�X\�����������O��l;B�`��I����ȃ�<? )!�O
<���WL<���n��������j��e���l��K*%����"�?�vE��-ϝw��W)��<ՙa5��Dv��."� ouQki��l���\�Y��r�lN{,H�� ��>W�9��hDǐ�Z��ς��ն?�}�����@#��8z,��=��|�MӬʗ��$ZR[[[�����j��5!�Į�$����A��8���������X�N�~��ҋ�7��)'E�� ]�Vg��N$ǩ6A������z�@���c���A>ȼ>Ii��Ժ��ϯ��b:�́��&v��N$t��67Jv�&NQE� �uAC	���E�c=�EF#�Xd�_�]A�V#�X� '>�� �L������Y4��V�T���G]$.�m��m�~@�te�-�.@�pM1���VQ.˝�/��#���|���z5�~ߚ$�D��� ���BͲG9���o-�����O����C$q��r]��b����&vyXK�|=���%(�=��tf�L;��~���,D,�g
b����^Ɨ�Z��j�����:���k:!n����|Q�z)Z��j:�h�&�p۬q������q��ͱ�s�G�~Ny��� L��˝���M���~�:n��YO�J�4��L�;���7J6�ˁK����8�m���a6I��1���p+n�0��ſ0�jPl�*�ݯ��������Я{�a��0Z�a�pf�|�7�f� wֲ�+K@.�$w�
�(r�)�(w+�C���f.�Ʌ9x-�IS�@�T�����N����.Z�}R�0�G���YP�b}k�3��1|g��&(����ZK14@�9ȹ����jN�/_���7C��t\�
s<tM:�EF�ٲ\P�z�`RF�1(�J��ڳ�/M��w%� ݿߟ��ڊ���׎A�X�� ���X]�[�!��=5ǿB+F�ƥ���/<x0 ���1
�4f��eV��u��R�K��ä;�W�q<A=�T�0��%���ُ(�m�5�e:Snbݕ�Z[��8d:.M��4s�f5�!,X����@Ec�������MOy�BGBc��:�*��tFIr�: ���{�4�6�[�(��p���Y9958e,�]���g�"�%z�[��?xFz2��\���6��S Z�W<��K�m��|t���a��A��'O�z�����~{ǩV]� �"���Y��o���â�H�\�����Nu:X!7BxuA�� ;s4�-\�Sv=��_S��Ys�b�"���4�"�х\��y��ZN[�\�.*�Ib�xs���<(F�ѷN��OT~Da��9M�W�v`s���2s���(vq�9�� j�h��(&���+�1y�j���M��A��]8[��_���jr]����3uW,�QC�������6Dzn�%��0��MS�0~Ѐ$_^/\�-tk���D��Y{/�`9q�QMh�	��XȠ�J��l�ᱧ&&~���#�)�a�Dc=���Q��+@���� Ʋ9Z�u*�u���|��� h�+0�?�3\:l������W��܈[k��A�*�_���KO��2څc�t#O�.�ZY}!%��	~����{�}cM��F9N�t|3P��x$�_xa�[D]�e��1=��o�j�xJq@����,�?��k����>H�-R`G'�A�!��W�k���N�h �k���:H�rM�"�k\���<)e��%D��u� 4�AcD�H��.bZp��mh}X�f�哉֔��-����>��1J��	Q�W�@�7���6�!����?���f��J���hU�Еv����	HX�D!<��٢�Ϣ�e��Бq:;��q�RFY�b#��;k�	'!g��e��e�������V��x]yl�#�S��}s}[i{��� �<�:�bu9��ym�^y��I>�3Q)�#��͵�
��K��3R@�qMg��l�l�����ΤZ���h	 �.�P�5����~}<���4~�	S�f�9��zgQy��1'.ue����,��Ki\����S���LZ^^~B��\$��&ϕmivnh"�]�{�[q�@L.�:Bwm�*�8 �GD|�7���,����M�'��[H�O��T�EKm�Y�w&8�c�UV+
�P�k;}�9�e)���Ʀ�;�^���m?� ڊ�����aY��$��t ?|O�Z�s�:� �Je������x�~.�r���t��� s�mgz$w֚�8u�nF��}
-�<��\�Y�<6�$K��+:$_R��cOb�A$�VD��)�3+�ET��`30���"Z�>g+�|����ZZh�o��{1�x~�n�������v"H�x<t�jP�ޤ������:1l�[+�P�}�^��"���� �j�A�4/��A�������$|�c=I�>J0D�3�.�p{
^�����S�1L�TYE��i�#�gb�-[R�eD��M�9��;�:�{�VS�IV�C�9*8\P��}+�뀑�N�S��K�bŠ�x��Qv[o��2R������}i_h���bd+y���ʰ�� ~|zzm�G���^P6�������AX}���k?�����;w���B�7-��:�y��y8x�G�~pF�Z�6�ak��r���v2N���~*�5����V\̃C���X��ͯ��,E���LL�-���C#��'g���e�7X�Mؔb�Id�p1���� (J`��1��֎��a
��=��@�SS}�x���������\ �^=_߿
�Lx�{򦃓҆�xOANT)�W:@R�����(����#C@D^Ow��T���zR������֫��[�Wx�P{hmk����"��Ɩ[a���ۼ��,���A��Mn�"Nx�4{'� ��'����Z�2V�?�wP�UR�*�)(**�v瞼l���dblL�M�����/�G� ����|�)��AIn�+�-M�r���A�2�&�:+�ev#d�5`�L #a��<�h��:��7F��2<�Z�m{���:H,�n���ֹ�'ݕF+��;�_����a�I�s�:�g��F��b5sLy��<y���	��T�h����[��A�����C�G ����M����.=E��5YQcXu&C��`�i���,���Z_���^�
��c��R5�������4NXx%���U(�"ҷ�՗ٌ6���B�5�ͼ��M��Oq\�3 ��D�m���9I���k������� 8U�z(���o��:�E����#h�ɤ������˙�l�P6�&d䦬2	�=� `CR<��9�]:�iײ�*�ַ�d�Y3����Lp8��r{.�\���0�R�����A�����$��Ar��� W�{��mQ�������5 ��ie�����uJ\��ݰZ�[}�siC��\����i���y�kZ��J��і�J�����M�l�T>�eC�-����~�� a_r�,�Q�`�^;��h��iy�>�5��N�0�tt��m�/��^|:�r�E��+'�15� �����ɵ���Ms���+��)I���*��	�Vt�<`p�o��󴑎/9w.3��jZ�"�X��~&�Yг���ϱ�V�l��J|�;׮�:��)-�ҝ�e���\[	cix�8��%.r0Ny-��Q� \���Z�ʬX8k5)�nJ:!S��yv_��A w���Ή�TR)���b���y$o0��a'@���$OnP�J�N�f�s2�����N�~����>��Za�	����yv�Ԯ��u�Q���f�:9T���%r����,�~gkE�w��EnuoY�����A_�r���:�o�`���\�4(^�(�Ao��͸�2C�b3����rx��Em4�O�k9U ��k�!�=���p&��R��@��:ֻRu�w�>�Kˣ����7���tF��2ݎ[$5����\ղ����z|TiR�dZ�nK�"�Jg�J��`Z����T(����4�V�W�v�߮��В�G�������:��[l��)X.�T��r_��`�l&����C�J��ҋ
�`0�~F��#A����E�#����ګ������ ��[+Y�	�|®�F�-��Ia����:]EC��ϟ?at�^煟���>�D;�v%Z�(�B;\��Q�q�j
���ޞ�_��k��B��P����'����mu�n�W�/&Į���W�GK}Y�\���&�T���^�A������W?A����o��8��m��^LX:<f��͏̵�G�����೑��\oS�PY����h�;��t�L/|�(���K+���γ���M�,6T��L��e��K'+3ׅ�'FF�y���s	<.)�1���E�@��K�8"��v�����7s�Չ�ouU�ˊ�+D���pi�u�o�Ξ�\h�����y�� ���5l{!��H�E+�L�{1�∐�Sy9!Ԕ�7GxB������\V��~?�5.��>��0���o�XZ�r�y��W�%4��z�?t^�E��y���룍�C�t���4�nsq��?(��(��@/��9�Jn����tF켎�c�Q��5E��K�8�WNV_� �L���ڐ�Lˍ�����Kr^QkX�AX�W`����������a�Vݾ�A֋ϖ�%��I7�a�l�ka
���"��yd��������j ���,��������x\y�m��(�G������wsg�7ޚ
/��B�h�g�����S:���%�d�8�n����2+^{�݄�`��p�F�[F��-Yޖc	��>#�lb;�q�>z5��$��b	��8MMM����L_�4<���	��E�u-,�;Q�Bj˂a����D' Y+,��q�%IY�����M]쀩.�R�B���S�i����Ъ0R�ښLv�s�} ͇#�0��g��><��.m�:*�t�p�ȑ6s�Eq��`�@��S4aa�i�꠯��陃��GPi� TO��ή�R3�	�P��e.��R�&�ڵ}	T�D�%����ȫ�]�Iu�mZU��O"R�D��:�
b���\#���>��T�\���9��Z�%���& ���ΡwR�F��s|�gUT�И��Ŕ� ���x���2�FY��qF ��s��Y�7�X��:dwfF�A*"J���ypn��t��-Z��� ��v��A�h�w��k.mIR���i�!0)��/ޓ���uO
XcU<���Hm�лb��oL}�kd2��)��H��)���W}4Rmb1���W�� U�#RL�����Z���GM=5�9�`�p���a+~��)��Fk>�_�Q�C�7K����RGǓ��
�"mB����,y��m�͔츢��[��磻����z�y��9���=�Y́���@-Խ�4S����-�w�����#��P�/�+bׄ�UQϳ|�#ZRrfԟN��-�bE��_{iX\�`k<���T�]�F�6h�F�k�n� �S��vyG�ȾYm�����Oj<����y�����PP��sp�9�.�ӥ�/���|�U��<��foz/ht���/��7њ���CR��ݻw؜_���~�G��&6N�~�,*�j��é�65k�{�۪iz��7�?�9�)��������w�� g�Ǻ�e}������v�({�"+��]���2ea4P����1��S\�@KK+ªQ��M� >ABR,.(�mN�򯐰�y�d<�[RpIHSyF�������C��@��͊��j7�CJAkt�����)��H�'>A�H�8Vp���U�t
�nk{�ݪH��^�cz�����4M6�C��M�ⴴ�ҥ��Ee,	%�ښ�e�0���f�*����NH��?��U���<h�پl���G�7!FN�(:$0ȸ��+�n���c&}����]��)�sW��r�4�}1e�<Q�6��m��ӿD|,b��7�Jh�\L�ly�w�G}�0t���2A�22P�s�c��B�Xg�		��~�΁&���O7�����?@�7aW�P'�����
�60��ݯ�S.�����Oa���?Tx�B	 f<~��0�N��Sm��� Ę��ZQ�����r@������AѕH���N����Ң��L/�rAM����JՐ2�=BoH:�|���@,�ά����)ڲ��l��mb�s#���20�"��7��5�����9ݙ�xi0����[���)0�Mi	��`���HW~e��5��+o�&Ӕ�����e�����cq���s$;��5��%�ɓ'7л5o�ۍ�rN�?V�n�@�M��T�q>��M�h+�؁Wb��?����a�񻉹�P�+t�,oC_�e4��x�:I�K*�U�|k��'!�*�4P<H�`G����m#��,�?;M����}kLn6M)N�1�^8f��+_7=�����򶲏�yg�ҾŹ�y;{�O��k�OS��U[g��C������6c?��g�~/;��3���Z�2�E�O�{��
�?���Y��-�L�zZb���t�/!!'.j��y�op�Vi����Q�?C�zu��{V�SGGQ�������"�*Z[[�1,M�8t3�W��(֔��:�~��LD_��&1y�9O־aId�q�Ӏ[��g瞦�H���s@������m,O��l�����~9%/O����<�U�x�e���YY�I4�wh�:�5�����A�n��B�s�S����  ����77g)��V���Uh�]ߺ�6T��TP�	}�������n���r�b��U��4��o�8�*�ӌ���	�������7Sn�d` o�/m�x��k��nc3?,̳ښ��$�����Z��(ּ��̶L��|[�3
���jT�����}rl�׏��O�U�nHS���	s�?+�n�������վz�OCC3�� "YR�ޟʥt>�x"��{dH����
Q�����'~�㇊� ���i�.=�f����񞌌LA� ���l4�StI���ʥ
�_uAl#���]������Q�R�}k�~�=,*j��>@oc�Ɖ�n�JK`���QF�&����H��>nQ�08��-��D����61>��P楠.B�[���Ѣb���ё�j+�NbR��=�N�%F�*�n�[��G=6u�N�~�����
���ϟ[�`H�#�m����"�/5�~1eE�+�7m���}wXx��������Z�v�g��?5~�f�`��|P�3~������\��neG�t�yڑ:wW�J����0�~�ܭ{eլ��1ɼI�sV8�L���I��M֤Mc�aYF�		���Moo�C5��Oq��Q#HiP؊N?���R��]��јm��V*%�E�\�Ĳ��UC�g)�k�b�=g>�޿��������`&��g��/>}�����s׾��SEk��'���^1|u����?$B�.s���E�K��ȩ:�#���!7�:5���=n������<c���z�����5Ȇ���U�Y)S�»�����V'�7\��?�@z������[�vܛ��B��[��@��W;#]K��F����~���O�9�-�̪_��kx*�7/��I�֣����+�G�Q���F;�[K�J��뿻n9

	�ׇ���������铓�\چ�$���/��jh���������������W�*�Ʋ>��KF9�s�s}~������8WE�e�ɗ��;(������h�Y�װ ����K
��(4gH__w4��}�C#[z�d>B8hPX�Ǐ_-a�14w0=��3��H$��z����G&�ꞈ�p-e�B��S%� {q�̚�Sbvi��EEZ����M�~��|�x���"j3�Z�fb�>;�u�`q�K'��;�B\�4���8�5pԭ_N��u@@�M]�*L{���v�3I��닾:�� ��]ˇ����C�o�;��#@�VSKB��Ȕ*Y��N �}�k���8�T������fRV�4M��l>r
�]����{�OF.[�T��'/KH(@Kv-[&�֨\Ty���֖�������@RɌ���JA�Scc�gA� ��L�>H� ;��|wB�������3})����Ҵ2ff��%���-Z���yi�������Ѿ��a���8B�#���ek�X�,�"x�Z.��{����"a�������S�P����`�{��d��Zjl�5�s�[3n��"|����ea&��DL�_� Wus��ľ�����]I%[�f�����
5�eg߿%V�5���*�J&IMѿ�h��Uz����=��1��.Pؓ@?��N������q�����)Bo�j�+�jIP�8/E0p�o�}�2*�{�y�^�B/O?V�{ԟP�$����\-�Ĩ�.p�1���+|Ys��1�����v����H��1{���P��_a.�����J�5�����3��90�{o�����/��%!86�v�c�U�u�)j�,��5Io��Fc�dn2�����(yyy���0��V*0�q�����@Iw��g�{t�=���n{����"�¸4���!�d!-H��a������U:��^V[;��������88<i/+pzdB-Y��޲!Jm�9�Y�D����´�
_�u���E'��WZ�bF�CB>�#��-,2 ��pPMAcN K 1���9a;���0�w�.��@��Q#����k�zH��&�����369�P$�Ø��Խ`Z߀7�����h�5N8ő�Cz�7zu���6݃�a�G��t�n$�˘Ï�;@`"?|8q�
����X�Gx��W#=3SE�0D��C
����:����,��kӑ��6#((���`}���1��н�$�$6!�P-������]����8y��?���]1����̑���&���^W6�v�L����ٽ0���K���+md�{
ǀ����c����G��'2	y�0�
���ۣ��.�����@�˳L x�N��S��&��$T�e�ȹ>zK����a���WU�hF�� �0�\`g�İ��fa�+Įo���%�2z�>��f�X���Y�4V[�����u��=���a=��z�>����������?��[�s���s�"�󃠑�,�>CCC�Y�h�o���MH�{����'���(��)kS�_���\{��i�Px50���Ԫׯ�?��P��3������K�+A���#���<+v�7Y�2D�������I�|O���R��h0���{��|��ӾG��Fȇ�p�k��D�ؤ�T�.�yz��C}�ز�4�:kR�!ԅI��'�}�3\����~�4���gdl�����R�0d w�Ő̾W���Ձ��^0�AWv[����������~tD7��
	�}RKG�Q0W���P�N\өg��4��k��X����@�-�P3+HH�7��O����R������I���S��d���SOa\(�v�,�d�#�r`�Ԥ+��5zŽ4���*����+��miZF��f���W���!_38<܈P��B}�� e�;��<s?Yj��\����s�`���0*�U}N�4(�w��_��z���O�zv�`�
��gk8��4�w�����{#�e1|թw>�F� #Ct�#X�..��Aк��=�K�l��SJ�;��B��d��?��F;���K@����Z�m�g*���	|�7�",yA��´`�2�����,#ZZy�+��2|O��'����a�e�M������D7��w�1�u?$���ѽ����fsJ�k5����Q`7�F�_Ԥ3S������oN+�������~2�5��Pi�n�e����P��q5�C��U�O,.��W{\7�a��&���Ƃ�����L�qg�7 ��Ӵ@9&���jO��Ͽ��R��\�A�7���h܅H�sg�n���wY~�{+�%��mgk����'-���_���	�WcMZ*���E�5$�Ȣ����w2X(�~�S��K̘@J �?�~=� 8��!�<�˰��8�~��)�yY�-ɤ'��}tjh{cF��d�P�{}߾}�.[Tw��մ�ӺL �K�]�x��U*�����_}�D���c�TV&�\�.:��������ޚ2����K�ʂ�u�!���� F�	���?��sY	�'�W��i;�kB|썏��RX�s5Lou�G�3���{�7s��(ۆ^\���	+������EA<�Ǯ�����
y4.����>�c����&�od1'}��,�-Z�_����e��1��f�qRc���@��J�!�_�����=��^����MpVV��� ˎ��0�	j��Ft������n�h%55����F�k:w���\� ;T�^}3�����%���2=����T��o >�)88x����SR�`b~�O���ph�� g����o	����a�{�6?�~JK��.�҆�"̗U ���_����Fg�!�BbRh�er�,���g�l�8*�93���7��
�)#j����~Rm�@x���S�а���Q�f�ϿYF�����d�524��%��Pt����o��6-�֡��AӦ��A��ou���K|��E�f~�J�et� �)<:������0t���������_%V�褀x���ƽ�bvxBe���/,�mJ�l�0�����3x�1���)��Aa�Z���$��e�[ܑ���@+&�uV�C�!{f�mҕ�i��,�>�2�ԇ8-Ȁ���N�U��ׇ�}K9��Z���?>��D������w�FAI�'Lg����z�P�G�N
Z����4N�?�$����~�/0T��0��V�h~��� ��3_r�ҕ��8?:��@ۜe?x���@7����}U��Gȯz�N���wXS��	MS�,���ҜS�e�y�Αͧ k�(�zH�>�9*�r������8 f.�����A��=�.���is���Q+��iᝥDUβ�~���G��O��,�{�n!s�
FB4�G#�Х��*ߥJ*�K��"*XHVI�zlBMK�l!��i�d��f��$���=�\��.[����з��rjs�� �$Щ<+$�S���&&�����!squ(��Ǐe��T22��!�����ĸ���!<L��2j@�����=�շ��˲��;J$Y�ӊa�Mb�)(((�i{�
 g�����m��(��&���Kv�q�[�;��v!������7���=�y�֐Gs���2�_�;�3I�}�P�G`-��/��,M�I�c��������k"�j���׸m��ik����&Z<�3{�^��q��,B���z[���9�C�$e񹗄��~��. �Ur�E�����|�߿	Y��7�X �y��b�e�I!o/}��R ���=����]����i������
��BF��>��6x�x��u�O�m�N3$�|u^2<��=sX&.��U��a3n$�����ђ�ɒ�չ��!f�ᑑqO�͏!\��di���>�?��m�vW�
0�p���^�s�8;�Pw�\��Pf5uDTC���c�2}ՏR�>��|s����"i���.<�S� �I�6a�~���۷�� ��	��c�c�.�H���i^8~���w��l91W��x��1�*"""����ћ�l�&&�Nq������m?�I�c��3z9�Sa����Q
��\'Zz������5XGa9��??��#SV�8�)tK�BJapܞ�;ey�7��.���?R>j��yN���6ַ��+Ao��d
P~�9h(J�f}�sX7=+���>u�4uY��a�/�C�tݚԙ�����M�Ͽ'�Zv�6j�diTD�
�frAu���ќ�ę����&𪡑�>Z�p�=�m� ���d~w�����p��a*W�U2��o��s�v���j\�eee�a�2��h؉`yz;핉��3��g����$���{�k!�%epV\�z�yk9�$A����ظA��,��ΐC`�����<���qe�Ԕ���Ҥ'�]�>0���U����"󏸃�|9��H.��jq{���S+�IHSU!D���e�
����!iu7m�Ey���j+K���$}��L>�5��{ݕ{F#/\����M�:�bX
$z�O��$��KC��Z;:��/�ڔ]穎�ݽL����x�Y���\**����_�d��w���i��D3ʨ1���G?����^��(	����j?Cq���7�}O�]���ʍ��?��Y����k[]%[����[<�]ٌ��$=6�Z�q��{V��<�h3~2�����q���fu�a�J??pD�}�:W�����|V��?u������A�T��#�1	r��ݿ�����d%+�ԓi�d�p����Fo/&�#�gÀ��lt���Ӌ��u�dC(�����������2-��Է�
��RN��A��.+}w�P����~����ő{k�ws//�W�<"*Q�5�*D���5��;v� �J�������K}[J���Do�ߔ�W�-w���8������:�^�c����ܽ;���{x8~���א�����J�U�ĸ��{=D(�fJ����]�xT��>h���]��6j���@fì���p��Om��������K������4��W�;_˂�b��KC@����[�ٙ�Y_krKӫ���p�����@�jc��	|�ʡa�N3=��9�ua�Н��P�����~e~?��USc�_���_J��c���Dl��W�q?�t�"�Ze�����|��g5���c:ۙ�W��Z�s]�\��69QE��:���$�b�O����͹�&����_��M9;��{ъރ�u�*�6�5<<�M�jU(��wM���?�!�|*M\-i���۹����=N��AEuC*T�<�Ql��
���xK"K��zc:g�'��ږK&1��[�dnI|�7����5�H"��t�2X��bR�f�Ұ��m���U6�O���c.� Wgt��*x�2!ҵ�^�7.Uf��ୢ[�+�,ᓑ�W���cX�ښ��N�r���R�~�+��,�帄HC�_Ev����M��\/�Y�8�ﳾ�&j{:�]͹���~��uur[�+%�F�E�ߝBR>}ji/^�����\�q��R+N9�����!ޠ;�5�ؚ-�-+�9~C�A���
�I�ܓG0;7�Q��R1�s��ُ;g�ip)E�uJ6]mU4�!��F1��BBj�Ɉ��lχ.����v!��"'!ܴ�mۏ�=/ޛ7q���~�l6�3����W
"�ĜA��,�LL��my�����d�-�0L�I����;�z;ܟ�����X�AT3�>�_1����Rcc˭�O��s�InI*�ԊF\'y<El�G'd���pr:��M��7��I�ses�\łH1�~54S�rv����ͦ\���7�d䗗�@ls�t���$NN�o�y��b&aɵB�Ah>^�T�-���n�-��gҕ�x��V�ϵ���n�ס�)۩^t�211������6M�?��;�OWV��u7�� x��(rDA��C��;��n|I��$Ρ���t	"%� �]������g���s�1�\{˝�m��9Ǝ������1�e�W���o�!iN^DuE��(.�6����5�M��>�M���Z��O��++`f�s�F�hƦ���|Μζ>�������]��2T0����m{&���/uԝ=�x�K=����%�g?�^0M�ʉl���\5���q�kR�o���F�1�@_N6���]�d�m y��S<��N�m�;;��ހ�^{�B����Mf��OT���3�F�O|)
��K�S	��`����x��B�y��ːcnf/-��nw�m<4Ռ��΂7���g�����T�}γ���[�[�:��Ӣd����rr	a~��u:�>h�<-c +m����d���J�򗄡|��ab���"�RA�_lY�Ue�N�P����6��EL�p�O�Ƶ�=˥�l@���� c��5�kw�%��Ҍ���|�6\,����9�9��Om�,6~./ݟ�}�P�b��n�%���Q�N��::��]��'z_��Jk���+��mvs��:���r�)�柟.
唗9&���{)�1�Qxc�|���^�V$�`3t��o���B�s��2☾�3[n��J�^�%Kܚ�����������G?�������Ù`:�W�m�n����T:d����A3y$]�.�p��%��@�_�����\�҅�WK�f,�8|W��0�W�zɹԆ�11�Է7����HX�Z]�M�
[�y���!��,�N���Y�V�띚J]2��?'ѭv��e�Ū��~M\�p �����a�ѷ�
O�G��2�9�U���H��PE�~�z�	4t��F80e��w`�`G�8 �>����6Zn���ȭ�����{�����(�Z{�wa����ԓ3)����*a9L�sAUT�v$��-,�z)[U&]���:�A�K%_ӉC8JĀ�G`CO~�z��fw���T5l6.l��}���3L6��.�����ِ�Y,��[.���-,�prqY�������j��f�����$�-J�����}f5�#t���Z�/RO^�Y�4�YĘ҄{қJ�6wPAB��S*_�*�Vº��Wy̗��S�p���GKŃuUUUGJ�#aC��A]�8.����q�O���ߘ,�þ�S�`�|<�����K	��h3X�
�4�*Nf�ğ"}g��P�	��C�M�P��G�6T�Bqџ?��8�_#E ���/��Mn��}��20��V�j�B� ���B���j����I֪��FƓR��Dx��	��-��ԭ���`��Y���SJ=2%�#�1��,7��E��p�^F�fq��R���{��~.�����\�$5U�*������[���>�Ϡ���b�[��

Խ�j�[ ,I�nJVVV�ާ###����l	z�ܟ���8`J�Se�BT��U,�T[����J;F�'_���Zir�K[�H-^R���*O��X#�ɇ�0�m?� $^���/�L8�ߴ�l����o�}������u5�rww���>�ÙFI��"F�	 @0�(�ä���7I�.{�*{yd�F�j�$��)cX#����g���_hT�)��s�>P��T�_]]����L��NNȂ��HK�7�j���L��t��p����O�D���b�3�;ct�/ Ϗ��9XXR���)('#à�,�(�ӧ�r�rsWZ�����w�����֤���;%�*��w��7���Q	#r�]Ի����r#�cM�it���[�wDkU��������
���o��.~Y�%�ga�w�{����D���X$�f]M ӌ�:F�ڙ�O�_[Z[9󃂂p����1Od��_ڝteeei�ݦ#×NH�v�:&�u̎�Ne=����1{��}������%W��!ԙ��B��cE*�iH����J�e�b-kՌ%�V5�	f���y�SO��
�s�%��#�!(Oe���@��W�'���V�8X~$�/{|hh8HeGф7�^t�һ���ـU�j�[d�_�ܡ$�S�'jϠ���_H�ʓ�!��_�U�?8�"*��07�11��o�i|/>�&��긝�Au���;܀&L$I��ܫҥ��;8+�4y��nA�������ZZU]����ӷ<���f�	����w�D���SϾB�w�z�~YIzO��{�7kƷ��{�}�p��P��mK�{����Ic9�rX�7��~	����RZ�Q� ��_Oh�_��)?X���&�y0ǀ�B�BP��{�M]� ��o۷��[�h�VG"����!O2�dA!'�� <�9}޻�_J#��s�w^3_�g�iH�@��5h�k7Ɣ�n ��$��{qy~���gy<�:�q�1|�K��c��(��#�tr\�H5ˬ�+����wu�
���b_;>�+�/�G?��S�.MޯbYe�$��-���B�?Ks�<Gk�O�����R-M�ڒ��|>�v�ᲪL�5�ս��%<�&k��4�Y�l�#%z�Rj�~y���`R��>���7��~p(�%۩[�y=#O�Bj��*%�حC�w��#����}�ͣ]F��/a-�
3�*�Bd�1�G�W�� h`��\<�RfÀ��ؑ�{�6��-ͽ7�����n�Pw�9�ac��]b� �b�.����$�Rmb�;�MT0�l+Xߐ���ɶ*pj��^Rv�&݀lE1$?ge����j�g���l<����{^�]uMY�;>ǰZ[W�2p�>��]xO�h"�nh���j����ದ����s�%�*d�! Ϭ�E%'*h��ɔ��mc�g�l�[�oh��KD ��\v����������BH�5�H���S�%`�B/�	��A����o1�L6<֌��M��U�(���E|S�o�+�"+�/;䍟��q��Kǌ��2���џ>I{oH���_�U1?���~��L��]����f�u{뽆��^9M� ������<��å Gq���pee���B[��IȮYX�����>����x�ߵMo0�?���\�Q��tNN���S�y�������zL\��2y�ӣ�=97dK����Yl��_�]��{���?��/���k���]��?��GE;;=g��&�����5�NLG�[�>��r��ߺ�z��O>��s>��7�bZ��06^��>y,���.�3Iӯ3��9�����8{�|��3xޢj���M��J��>�*"���M�k�D���tu�+4��ĭj�8?K��{�\�?W���sb9T��ȷ�ڊ{�SL.���1H�q*n�r�{0\L�FϿ��x���H:X蜧5��-M��7���,�(�{Q|���.���j��2Ϩ�P+&��60B��i��u`b��c��k���f���=m2csԊh�6.S
$���:����h��hE0��jW���]ݻrF��U�΄��r��'ÃTƧ!��/�o��\�J��G�EmV��|��zGz��~���mJ	�u%�Y����{df�5bV�(nt��~3���0���^��5�6i�g���O99��\�;"�O&Y5Ruoe����G��<m\,� ��Q'���4��K�g�̗�?���%�5����w�e�筜�H������+oKM����_�d �Eo ����}��Ӌ/!��G�ss�ܩSܻU���n�1VvV�x�Cjr!C��g��OJ`��8��ṬW%?>z�<$;�Q���wy^�i����ZiQ��S�;�SQJo��C��Yhx�!���|��6v���R�5�p�b*��4��(԰�[�*�G�������+B���5�Js�y�ai��Q΁M�Nv� ���W���cuj��!|�o�IV��h�@��ϻwğqf��\���wF:n����I��?�%]d��02�n���T[koJ3Ś#����׫���#f�+�#iEX�w�\�u�L�2��h�`fPᨨ�j�f�����|�^�j�K�k�lr�#��X�\퓉�OG'��ad?�7�8O�G�xPO̼P��f>�J�_�{��;!���S����ɤ��65Ӽ8�Չ����O/+v��H�9�J�QŃ�����}9F.?��g�����ԛ�(���lֽR5ë��wP�%�;S��h���)z����U��-SKͺ�s�����L�-Ug*O��.��f�v��.��hk��]�e)����rܝ�>��/ᗹµ�Nᮞz��U�l^��d��O��/[�TRQ�e���廻����1��������qE���Ń�R�UϷ�f*S��/&#ɐp�hg��F72�>H�3��^�n(_��4����-��5��튛:��"c��tj=%la�ngt�͍�e�ܜHg	d� ou�*��c�㋯�?0�"N�mJ],^-:Ӷ!Y H��1P���tY��b���.��j(g����_�
��7i�N������ ���zY�x�L��x��z�ق�2��vj&��?]�NAw��3n�<a8�����`����D��-S��N�����歔B\"�ѯ�#O+����i����ޕ5������co�W���l�$q6��!a���*ܕR�lq>z�Z�`����W�y��Ʊ��/#�皩|Q�!�*��z���4#R���+�I��W�l����\Xݍ.}�m�N����Dc�11+k��ڒ
���F$��a��3}�������<g[=��[�[���f��8�B�~D<���V{�����ڧ�8H��zE�+��N��TF��RQ�ˠd����m����l�k�j��m��H����RaE�2�����P�'�_`��JGwM�Q�<z��`Y��:з#	�[����'.�j�����J�.�e*�O���;e�����?��W�F �	�������g�m��LgNr*jr�D훱#�7b�m���U�J�P�����
����x3~q����")i`� A1��ڇ?_������{n���
��"%�F��`��r��M�(�om��'݋eg}�2c�\���h��T��ŗ�'h��#t/*)�:'U�Y/?����nE������=��
��{.N���鳰�RE��R�
�Dm���e��l���ꤻJ/qC���;y���"�,m�N���t��^̇i��|'�<�����';q�5���|2�R��iO��+��'IJӌ��㒎����j>f}gs$�jt==13��r��ۄ�a��:�nb8iC��~��"f�f����z�__A��u�������K�A��I�#�S�tQ�?��%h��Wq=b����):Ґ��!H����fQ�����K�=Z=�椄O|�TY>�6��[�j��o�<��)������3f/A#s�G%�~R>Em�I���c^F�5��~��~�1Z�$�],��
Z�;\��*����p���0�2%����|�W��)K����[���5ϵ3��]ڣŮ�<�=ާ�K�djU\ѝ�8S��e�ƍ�Q6
��N�����+c�X�����G�٨��Kw��[r�KǑL�H�X�ӿٍ�����S���0��^y[3ƙ����
��-t��Nr��N�QJYr�K�q��''�j=�`��BV���j۔�,a�Z��ΒA����_5">�>�g�����w\���{�b]�t�c�T�Z�4����[�)f��o?��*��C|T�O/.y�D��S"�2��=�"F��?�]]]1+^^R{��CԦ��AN�ƶnQ��D����w�H��T�d�&�0�X��$*%M<\�ؽ��ߤ񄣩k���z7o���N�C� O��A�9A,�����6'2�ڽ0������V��>҇��l�7�̋|���-�~�,�q�Dē�"_u\�i�IR��.��K3��0|F��+*��I���j�j�N�f>=�]�'w#[Z�||�Q�6�$������t+��ry��u��Ϟ{���f�������g�)�D6<�?4IG�W,*VF��/�{���%��B��K�����8;��� mA�����p�s��ڧ.f
��8���ߩ����}��㮖��"!�9�}��9��c���;a��v{]s{�2��\Eו��<<��^.F��L��Q�v/��pm������)�Һ�oE�A٤z8<��6ˬ����Ϟy���t��dNԚe�Z����f��H�����7?�sT�Ȝ*�X�a��QZw�g���.<�`�{'O�~�lIE}.�6���\�ڗ�7I޿���Nå7ǌ�ީ+�-��l2�8#�k:��&���cb�!7Y��t������"��=�Y!8~�,����V�=����L���*�Y��|@oY������#�:��e{>S%!!���Bp�&�%s����`^˿x JQ��Ό�<:C~�`cHBD�;d4P��[{���F^bi�p~Z6Y��f���ί���]�;��� ������2���_�$��h�K���g<����K�����s�wh��l�W�%�ݠ��ɣ�f��q�+m��Am��,�sɡ�OMl�~̍��V�,^�(���sj��\݆'�G!���k��
e~���E��5�!+���" Aw>�MH��K�n#�X��,�̏�k�$Y/nx=<?��&mup������Oԝ�*��;y�wmn�6y<�!��k/Y}P[��Q���HAq�\�l������s�x�|`���)"�j�f<w3SV�i�WB�"*K�=�5�R�&e��W������ז�h��o���*��Elê�E`�.Se�A{�ŞPK>�����H��9
�P�禃xL�V̾��҇/���G��-�`?ߧ	�صR����ǅ��H�T G�:��e"*�S,Ke|��rZ�*2r���$��-a�mi#�o�������gA����m8kr��-��;;*���@�֛y9��BB��Q�M�`���"���&X�)�����#��_�W�	D(l7��t�J���QO&\����g��m������~L���zD�ʰ�S�b;\��Z��A��^���©��,�Y�~�wQK-�8YW���L�ȋ�H���T��A�ʠw�d�����UF.�`�=3bsuk͑Z��C��.��*�<ڵ���f��sq����	e�"��˗�J�EJ-��wM[���e��*}�t~d)��M�틭dk��_��L����^rY�6�@�	��i�3�������wm�c���TgV@�>W��+�L�i4��HPc@4����)��c�kO{�ц���'��6j�b�7@�2<��#[Zvc�J�^����|�x|CJ��k�F��J�<hCv���b����2c�y*+�R�Te�Zu�/��������e�	�]� ����-�XE�N}��9Q^kK�2R��������8���e6kr���#�x�Z�e��:f(%!1�q��!CI4�ϢS����s%^�k��;7
z�x��þ5�d|c�cnڥU���T��/?���4�g��J�-l6h���q/0��/Š���t8�@����� ]=ɗ+&��g��a�8<���rMZ]{�CƩ�M�C4\��eo%�C�v�}2���N�W豭��[��EJ-�ڧt�>�3����)~�W�/yӷ�j�zԪ�D��|��)?�u����@763����hM��Yn�Q����"�J�����>T���N�-&��f��Cl�.���`�7G�	����Am�8@��~E��򂈏.�:a��PtYą����<�N�.�\�ȟ�,X��"6̭�*��S��s��;ka|�rc��3wrV���'�/l�6_ L��ܡ6�K�C;�p^IvG>�����D�҅�Փ��o
F���[���#滻����M;��Jv�I�II4豵�����é;���L��<�6�j�.���B�D�+)m|ٟ�0E��2�q;��ӷv�6ؕO	���\|��v AN�h^`�F���'^����Й��#Ú��>g���![[���(�[Znu��+#�Y���)Aov6�Rb8?4B��Okۈo4���z8�<��[>�`��XsmJrep}��8����8�t�&
�ب��՞�z�T��|�}��m>���Y�����v����I�h�����m�]��5K
���Mke���LjIE'3Br���[��{`�lV�us��&w'<��7'��D��嚎G\�T�:;w;�vF���
y�$U.a�Ѧx�@1F��$�R��Л�ȏ[�F�H,sC��@�?0\��/>D�}w�?�[�B[-�}��ӫ}�6�!��_y��h��3�s/����Z`�z���T�x0��������ՅŭJ���e*����M�v>�8l���.`�,{F�5�u��=<.���̽G���e�2����j�nmvv��-��&B?���VJV�5�4c}p�xc秸[��n��9�XZΚ��_Z��?<~_e�K��`+``�uijp&�	(l{L�q�U5[� �.�΃	���rO�M�_\�~N�&��|�*p�ڝT��c#�0Ե�.6�$����ϑ�|�[3)��ѓ�؛�j�X�/�J-ژ3+kF�9�U*��X9�k/eͲ�ep�^��qO���7�Xq�	S�J�y�����K����E��>�c��C(NS��5�n+�l�����o�g�^2BM41��K��}�lԽ�s��d����]oV� �{Ցb����HbYd�5W(0��E���o� ��EW�s�X�״��%�������2�O�����7��=���95e�㕐�=�� �eK��/99��n��8m�)�If��N~4�$��k��c6���;���ȸ^~��2�p������ri���ؘ�MSD��k�7#����!�QK�G���i/+^�����1�T&/���60Q5�ܗ׭���(M;�e�8��q��/l��"S�X��~����ꗢ`!b�u.�1gm�wa@�WOU��N�Lg>?��a�Ā �!�i�|����n���{���\��פ�@k��uJ��~�"�G2�g.� ��k�<O� i0�n}��n:�����g�Y6�1/D'a&��LL4���m!ŧTc#"��5?�s��8�s�;s�hGp%K�
�h�3��"���1XQ�T�����S���\�i���*!ϴZ�¡�u���JY�RlT�V�>�yy`$�r+�o�!ߔϐ���F�	�p�N3��h��8/(B�JLr���Lz {M7��s�c0�rz:�aLUK���ř�_�x��H�3ej��G(:Xɧ=E�)��y^�}�2��'�>��T[[o�Ivc�3):{UVN�U�ߥdһw���)'ڄ����N�Łn�_)~@���L!uJP��XU�Y��+��������.B�+9��{+�(����K]��1�{��p3�[��f�>7M�Z���:��FW��Hz���)i�Q!��^�v�^�l5@�m��NʷrE��g�Zb��t8�n�|2O3�ME�zX?�H.t$�"��eFv�ï:Pz�ޛ�?��݌�o��xj�"#�p)K�S-2��4h޻YY����#�ՙ�]���c_����n�SD�9���l�hU���Dp *p�b	�},X����M����q��ַ����&N�i�Y�Ԣ����KU�M��7����dQ�o����y�#�@��|��"n+�#S��܇�jwڃ�s�4*�o���1�L�xe��%�Y��c�a�|��t"14��&���)��\�$oBR'K!��Ҳ_���j�ir�~Y��\�3A�Z��'��`^�iAl�I鎫)���Q?+��B��=<!�H��Pl���m���x��4�E�J�:���s'�bA�W�%Ӷ=�4Y����|���C��r��2n�Լ3�i��d�US/�L��6�)�7�W��f�ݺ��i�A��Y�&H������̡��~F`�d
��M�B#ءbí�|��S8��X�F���P�z4�e�~��;�����Ƹ�Vqd:���J���7���v"�EyH7~�OH%]�������t���A��'э2�sp��9(�Z���a�OP�`�jO�$���o���e�a
+;��V�x��/i1-B�f��ì���#�����3��y�W���P`�^�m{�'��g����:�V�i��?��wS׉.q5e��n����3�r
&����:�f~5""GO�~�����>��߂TZ�BR�c���.�v�4��1�u��+��T }��7MSwܤ�4�l�����8;"��
�e��@�TPAF�;�7�--��ȭ�����`��@��;��ݦ�f�K�5�+�5@A�x�$4�\��e9�6N��]]�A�}� Sō��W�0?ȃg�\r/��~�S�a�#+��O��>y2�¦@s�������a��k&T�
����D���р�\����;Al��mY\L���
Ǎ�9�>�V�L���C����*�Rg*��OWq�b��WVV���Q@N�1p�\��wp�+z�[)$>���˂)�l6�m�*c��iԒM_BN���3|y��&#~�M�ɞO�ȿ]��ߕ}��s8�<-�@�YY��ɥ�hk<�j[&b_k�{=vt������m�;jH�֥ �V����He����J4WW.� ��$�X��.P��	�����S�óa�ז'��ǿ�F #�xX�g;�ΐ�H� /Is�)P�)޿��9R�u�YФ�����PS�a�>�M
��f��~���_�nr:}ڼ6�D1�V��?8H�BW�jT�S8$	*�ߪ�㭗��S���V�i������lW�����i9���I&�S~&�LMR�戎3��ځ1G|u�:}|8���Uz�6^b��{�	.��f$�S����(��P�IÁ@5��r_�|�؜�L~H�����C�/�ΤDEN�gb�6�^Iч�O�+��[=,�;���@��y�?̚t���h�¿���4���j��R��R?���t��Q^���G�<ZZ��o�9=g�THu��6~Hg(�\����+c�N'�Q�@�M:(��y���v^?�IO*��V��44%&�ؙ�U�0��M��	��0f�Y�������z��� ��)�f��KO��^	Rxﴌ����H �8�AҚ-���iV�.�7�b0��[P�ٽB�ޯ'�rwE=/*I(V�S_ñw�����:�_��0Т��������.� ���i+�\���ɞ/F������L�C�d�j|&��AO��q%Of�,ٽO&�YM���>�&���'��"=ݯ=H�A܀�������S��&;��b���'&�����c)��<��j6
��� �¯L����빿��}*p@���t��T�B{��<��9g�} V���cmZ[��[9�̋���抬�)Qc������RP+"�T0��p=��R+dv��o����]��4�I-���S��"
��:Q��+e���%@��} &Ӊ�WL�X�����I�1>1T��]맅R5�J;��]�'�]��$^Y��-��{8G��
�R;�@f��|N��[ŵz�h�.2�*�Q�'�� ;Q��}Zi��ct�lh���������d/��[�����Ӯb�pܹi�d�iZx�g�­F��'��M'�6EW)U���W�U٘�k�x��.���9L���b"�*�v3�h����7p	���M�� �q���vnTi@�����x��a`��]Q����,f��;H�����~/>(z��ԝ[&�I����z:Y��C_~�=�]ST#��y���E�"���Ư :v�H��
��]-�?1p������`P�e��������5V�Qx_7O�V��t��6U���#\]�+}4跆|E�Q����D�7-�W2�Y�)Pꠜ��"�q��H5q�E�4<��6�U Bp dp��`���z�O�s5��+�y�dM-Ǉ���޽�Mc��a
��s� ���t�M�N�����GNT 	S�(:�=���x��ã6��ZX��J��.B��R}Bߘ;�Cf�נ=0��2�F��K~�%&pA��:���./��ǃ�M�r����H5&��;���|?��$��di��2��%����4��B���}��wp����0��o)z��4e��C���Z<G�$�+��u���#r���"����B��� ���n8��;�?]P[�g��A�b	�<�chH��#�@g[��v�FN��5�m����S5|ń8^��m�1ߤB�l���uPmA\��<x��O���H�|��
�'����)��)����3&�w��X��n��j�7���_�"�Dl�A��[�x�5���T��0i������0��}�1�E�k�Yو::�|.�*6�y҂EGX�����{��FA
����&�brJlH����]=��q'����SU ']� �Y65c�JB�4?�^C¡=�c?{�=�Ql2,@�I<�]a����	n��ۅ�5���L���a��٠�<��{���{���`��_��Af_���d<��L�][w�pbU�#N���W������"�<�7���������CI�s' ��'s��C͉?�?�ݨP�uk5�U
���՟�BC��\ 7�4q.+�NIm�u����ŕ����{B��3R��N��DH��6��H|�^�rmW��G�Yj|��os�<���|i}�IA����ڀj�7����ͬ>��*a��[C 0;������2����<�b�w��M�Vissa�۾���W�'����/캳�Q�	�Ǥp�3�@ܭ�ʝ-f�qݺZ���X��
��yy�2�nY��a³�Eާ�6���x�:�=�Y`}�R˸(��H�?�#�yQ:g�d�t�
bю����}�ɢM��3�A��K��>p+suUi�����o���tu��Ia%��R���o�~�[���)Ā��`;'��Ӊ�O�I���E��+��3�����B�̔����~ǣ���s9m1s(Օ� �`�3�.�x:�mA)���K�'�礭�����e«���-�4�3)�b�{���I�e��h19��I�m�^q�p~p�u
(�㨔��(4i!���I�%h�3�c��J�~�ZV� �����)�RRl:s�����!�����U-����Bx���Xz������rP.�OaP��Ƃ��L�r>�j>Xdd��EW9-K� �\�<���kt�)���=]�s[�s[H20��Ee�l��Ѭ���\!�����Ff���!���_��@���6c_[15$	N���P�$Ӄ}�=.�V���+��
w�2*����3����J��<��ہ]��S�����F�(���Z�^�8B�[kx��8+�}c#z�>�i߫zG��f4Dj��:��Y �F�$�4c��E����`��M8�Ϧ��ӓ�&�Wd^��wc�K�mz����_u�JE_Wa��@� �:_,0��+�;�$ g��~Ē�qg���)W�I�F������K4��R.V,����=�2A��/�2XP���P�-�Spciio6W>$����g8])��W�|?o^�I�NPUe�K�Lo�+��{fi%�{�M(Pq�# Ձ�|�XU�%}�;dvpH��*�V~h�7M��������b&]��?b�Y�l���+e���֊������D_�@��� �gކiڜ�ugȷj�lP���a��#�+���y`��'�n59x/�r='0贈-��65Tod ���q�Sn�w��>2?�eWCa������	 $�~��������q �G��ą���ShU5փK�������Fm
qxEl�	�=.Q�Գ�<Цv4��
x��DD���"�wDT�j�\614�4�%�-�xـ����o���F)������@�C���rv4���#+6p[��{����B�\s��B��6������瑵z*���!ؚUl:6�	�JR\r/KZi48�F``��@$�A�oߝ��"�L�������'<1!��Z��z�ꪘ�gM��r�\ݩ=iQ��e1�G�k�ż�ܤ�����W��V��ښ�{�ZC�O9r)d�I����!!���4X����ϊMK�l������D�
��+:�����C�t��a��?�|3 }��#y�~�ԅ��t��FӞ�0���
ɶ��ŋ3ڲnx�l������1������3x1�N�=��ʕŹ�jk�.��Ȼ����r��eB�1U�W�bT�\K����o���AP��	{�O�Pj ��)�+SWA�R���n:Flƺ��%�%l
ؽ��p	�Z����	�8V���gm�!Y��U������>E�Ĭ� ���w�d��w\��[����p�����	������=�y�]h���Ǿ�4�8]$�_�QdtU	��
O��t6���wEb��u�t�U%� ��5vҢ-���^g�͢м�HS� �E��}��k.���ѐ�+p�b��J
�9C�(� @���g`&czjR'�LN�1B��,�E��T���e�f3Y	t����A+�6��r�	I$,�yM,߄�~\����/)v&iNP�o>|G)I:�8�W�;���l���1�&�����	���$��)��e��|gF��&M{� �
�N�U��$��uq�5죂��)�$?��m��*{�?�}p-�	���mi�R�λL�"����[��u��BҜ��j-�*Z�C��9��O ��^���ҙ���͎�s�f�/�|^�fs��
�.n���I�G���Y�H?P8�F"3�B�)�|Bl��wӪ������2t`�ѡ���BW��bB�058�M{��U��T}�s /�m�Y���I�Ku��Kv��$�����u:2���>���ݟ|�Ru�(cO��$°
�q5���[_��ʙ�)Wp��`B�B-L���ݍ/��D
A�F�u�gF�Mc|�
���壪>��%��@�	,�ن�P�����u��Ҟ�Vm�����0�oʛP���X�e:��v������a���э��ա��KBt1��Ho�}G�jP�Tw`�mp�s���G�-���^{:�� _@�G?�7@���C���G^<B�n_(`d3^���6�i��H�έsg��9����hV5�t���Z�e�
c��˻��{�чqQǵ�6�I	���p��Ո;w���b;�0 |�ӂ���k�:�TW"���E����A�s8��L�4�<E��k��{�t��/�' �߂�:��z�_`tݢ��8-�Q[���?�c$��ϵ�⺗��i�b7�� .�K�� g#� �y�Q�x�Åw����H�������*|�&uu5%��.rc,(�|���@�ҕ��/��%Pp�^�Ӕ��~$L:n=;��R@>�hr��%���ݨ#W�{
��R�(�P�G!P�;��0���uA���?��������7��jW����0[=J��7rϤ�	Je����[���y�����IR����iCw6o��P�3���qE�˛K,(XK��0�x��a�$�=�6��=[�'���AH ���5��}}K"�bpO�j.
E��"-�u�\�Y����httKبF��NH%-�:P:�C�}cH�0������*�xλ�;y�9ti�����ғml�j� e����8T�No@�~����pTtt�d�㮂i�b��ex������O!��]�auwֽ4���Z+��~����|��k��G0�P4�87��Ώ�֜�u{���B������.�
�,v�q�d'����2�u�D�^̟�W����[�������@�ش�\�5.{t������	6KEd�2�7��l��w�G�fL����?��5��&y���~�5W�*�oH(6٣I6J]���+*��<�޾�{��j0���=\1� ��֐�-�L]^.��0q\|��M\���4��A
$B:�.�yܱ�R�6�ՠ�x&��'ܧSGv@�5<B#���<u0�ø��Yj;�텈E��[�c0ٯ$>�u���3��p���eR_#T��� oHa<�kZX�q��0��aw�nZ^8��U#�ɝ/�9��홨���DJ�D���gʱ"_7�� "B\K�GG^�Lz#:�i
�|'GV�Uc��@�DJ:5����'׋T _-:��	�N����n�$��8���������߄������ ]l��ڑ���}�s���+��h �RF\U�ʳO�`C��KP(p�)~��;�e�3�_HX|�p�? C��W[�C�9i�6^�擇pb�=⓿����d�ܼf��u�I� �C�_�i�׼��~n5��;�g�A ���j��S�@ee��城Q�T�9y��0�.���\���"�_����C�\�Ύ�i$5���Dp�4�]Z{�c_17K�_!����;^'M:H?8��0���j���mZ��w1&�?�t�Xަ�<�����m���c��x3�RT��8�f�\5�WKc�m�U��}/ ��p�T���s�	�'2�<��<���]d�Wu�.��p�=�E�_�M�WVV�X����k5pD:0�l܈�jx�6|}��UHBby}��E��O�@��.��}rߗ���m:�1[{��-��0��~�L��%f6�w[Olĺ��y��`ii� �G!=�ԋ�hJ�����'T�բ��J�ӭ/�x�{�wSm��6.�z�\S}�6�֠��vͺ��a�8�+10Z����ԇί@o��x�;P*~j�,����ձ��~�ĕ�aA��'��䭙�	�%��U���0j8��;s�_�@��wtY�Q(W����;Q���_�n�ĪL�����*�Q'�ɰ�zaafNg�_���0����q�4`�(�C(BSWν����ltX��,V'��?]l[ւ)q���B�Q�\����Z��E����p��<�����0���&:wO0�)��
����A�ۖz�I+���`�7ʡ�<\ΖAn���| ������񥿮)V���F?s4�c���U��d�����W�y�#6���`�4G����re�Q��VZ��1ؚ���[�Su��q�J��/S[�T��tj�t�R�Z��ж�����:����I�~'[w��L悔@�5��W�RvYw}X5aC~�r����Z���a��1��\�m��6��"����Jn�h���	s���q��z�+'�%XMو�|;鄯��]>�U4��Ce+�1�4�o1��L�ϱ�N�s�r��T������]�B�}�n�S�#.RL1V8+��p+�1�k�f�F,8�OFT��>����i�7�����\����V||@�Z�߁#���U�H�����2���KV����"�{�dfs�%J";�ڄ�E������ڄ��>�����?��~��y=��}ν����� �ISK��V���H;�	� j�:Cn&�[�9�4Z�~�v��z���jj5%2�8��k(�Y	��������zz����cEr����/n}%!��q�鍽�ߏJ�����IIB�c�-��S� ���Y�bڳ���J��!�{��!�n��D;4��q���~�j������U\4K������GO�ƛCC ���p�"��9��p!���	<���"��9�Q30L�� M�i_�*d���@���|e����5]�o
������m�3�.f�]$󔃠����tLڎ:UY���j@W�i	;m�������A�J�qZ��0����:��4�Ӷ�B�c��#2' �@�$_��a	����b���q=M���Y��<g��l�Vh:�j�U�찏��=�K2�ܡ50g-��9�8�}g'ͫҰ���-��s�oū�� �6VLW8�;�03�i��L�*�UV��pPm{�/�"c>�c�:5��X��	U�Զ����K�9�tϛ�P=-A��u�v�"�x�l�R��e���2����% /7_�V A���Ŝk++OQ��#g_��3�J	�b/��Ԭ��������	���9���8��00^���sT:���.�H���F���w�bP[Y%�ccg ��/39n�i����4QV7Z�%f|�9,-��ق3��oP�����.�TV��*xW�z��� �OA? ^����ҵOA��Z�Ȉ%���֨q0���F1J}$c8���^�%?0i�������ˆ����{=az��1P6\`(�o�X���9	��9��ǻnn�2�p�h�tyLh!�?cM��^��v<C���R��$d�'ۅ*kt$�E.����/WO��W���O_q"=��ՌJV�w��L�0X����L_GqN�~��p����3�P;.wHqs�5��.��4�n�+#Z�.���V�6��o���;�u�y������}�C���d2��R�g�B���/-b�蟏�k%����aG�ĺ��dK�Ԁ���"�{��.���j*�y\�߂�싘<�k���ub5WY�1{�+F��B�ི�h�x`mE�W��0�'1��f:�����j�lw�U��竫�G�vo�q��j2����B0>�<��}��٘���!�k˻��m�>|�/Nž�g�>��<�۽L
_��
%�<�r�9P�P���/1�	.#��D}ۯ�>n�4�@�\/m<��'��֛��H��{�����f�
n85�T���Fʶ5�qѭ�3�_N3x1��u��4�1� Wv�x{��X�m������%8�u�}@������{j�&Ӧ��)�6d��+8�Yc^O�ՐǴw '�����{����<k��g��	<# �=�dR�?���lKYݺeM��=1��Z6Jxʑ8�����ϳ^��	Li��r�����xr�De@���Q۪��
�󘲴���1��"�7ӻ$�����j�� YU�@��Z�-�<}X2q.�3����wfړSE�:J{�����	���_ ��;���&7E30N��z:"w��,O�20��F-�����!�rT���<p8<�o����P��a�`��M�b��NhW�l{��F��SGY��=��f�%W�X�w!| �o��,Fd�Ш�4�f\e�T�Klp�UԼz��;.u��bd|�5?J��љ���zO�Or�M����W�p{��X�rN��T9/9���}@�O�w�7f\q�W<��o嬄�d�R$=�nk�״�k]/��������^'�ф�j��"��2>Q��m\�k��^��Ɖ�"��S�
XA�/.X��h�q��W���kL	^2���	�UBY������v��׋_o���DJȋ!���F�W�l���i�B�wN�x��pw����{��ޗ�\Y&e�m��b�G);�|�2��N�!�qv��Ef�5<�,F�i8!�PDن�&mB:}Ƶ�巉�,�߀^���M�[2T�@ _fMx+6	B�R
���<q�;x��������l�O\������9��Q�!�|����V(e�d��w���ۀ�'��"s!���Q��=�*ן��˷�@''e���'��M�����Đ��ݙ�Q�7؟U��n���fY\T��ZE�������u�tc�r՛�̺Mm0�l�Ŏ�V�t�5�����-����ηv���2�w]�k]�3�l������ダ�	�i���D�v�쪶ݐ�ʸو�xU�o�[�^�f�ιJk�����`�Q�h��z��t��k���,0
�1�Dݴ�NkNX�&Z�Ԥ8)��M�2����.Em��Ѻ0$~���~����8�N��n���
?�.B��jnfӅ��>ͨG
O9��p�	���p�t��b��9a"L�E�����OEQ?o>S�.�t�.������'n�nG%<� 鬽U�9�]�Z 'g��y����	7$+�:]�JjF���'�J�Z���d��4a
��H�����L�� �a�P�	A.�E���=O=�qDE���sr��t}Y���ǡ�g�M,�o>����̾�:���3E�e�FWUłfM_U�g���p�����θˇ�+uv�Ѐ���m�����n�'�2�]�"�Niek�@�Yx�]�.�wd��vEU��OW{ �����\UeE���e��OQV��#2{� *X�~8�Km�����
bG�������/�I�B�'#���2��d�nNn,����!Mu����\��f�����B��;�ڂNE���߃�$�������ύ��3c��s��@��Nh#83'D�Ǣ�y� �Ju��ʪ<��0�j������{�@�,�K&���e\��,F���"���3�z5�а^kAaj�.�:㞇�VFb���kYM~���\v�=�O��$
)n,g��Y�#�?$�y��93�)M��~�<N�,,ﰿ�/+yp�Y�?�e�dp�}O��_�m<��'�KC��;�RO��0ϑ�0�ww��PBtmB2` h�9��r֑n��=��Eh7�iI�^�I&ZXݿ�hK_��}N��@D���W�! ���뫗�	M^~�Y�u��s��W��$7�Xt(T)��9ձ�23��v�q�T�
���Ӓʶ���5A��7��3�8зܝ{��J��?0a���.|!&ƚ����������.�wR��p|�v��g6�1�1��ZN������8�����ߟ1�s��x�˄��Ȟ\'��jAd/��6uc��Ci�5֓������;F�R��]�������zsq�?��N!���RW/§��p���c������6��y�L�n��H.�������w�j2W��f�&��-;��ÁB�.x]&�����ٵ���In���v�֧)�64�}��s�t4Afb'������Q�d`F�J�z�VQ��a9��?xl����75Z�w�����r2��`����{�d2E��zxܖ;K�F|�ߠ�_���,Je�W!/W�V�za�BAHo�L�%���|y��I��meĽ_�Q�"[f�~��pL���厮�w)G~���h�U?�8yʛ��"Sc���7D���#Z�[D^(?.q�X�e��u�Q�g��
�TF�\�m>�,|�:|�q[u���r�����hsr�!-m�7���(��W�94n;�~��-b��p	Z(bk��n��LY�
�`�a��R}�I�xU�~88�[;O�"���F���l�w(���]x�i��e�yr�&���L���P� u筚[�f�w�.F�����`e0��� jI�1�N���̑U�D���S@�9H1'lT@q�KR��Q�����u�}rk�4�Q�,D��ۤ���=��#/�$�l�`�|	����i���ջ0�e�=��.u�ka�*19�z^0lM�ת�N��-l�ڦ�����?\�9��5<������O�N=� ���I3�k�Т|�2�=
3��VK��(Z�O/NS]��=^�S�i}�z�& ��v�����HsOU��?>x-c�0Z�>g���K� 7�D�(6��a��+ĸ��B4#.�4=��v3i��%BTf�-� _��-����YÐܫu�0u�m}R��q^+�B��E�7�e�W���a�(_>��WRX�X7���o6�&��,�9^jI�2»I;oF+�E�۶&��3��%������>~�qK��,��lU�ǯ�VǂB�n��⛒�r�5o��L���Q5�	A����s>D��| ��-�?�23uͅ�2=�"����W��s*����p/xWj��B=)�)��Ӧ/�m"ӝP�&.� UW��H��z���}xO*$��[�4���1N6]:R�4�y��ͫ�@0�m]u������N(#'�W��5���t��]��l�V:�,�b��� ��TO��̽,�Qp5kǆpz_��:��
�Q��7�aN��y����Kn"ĨՐ��5�v��G��^	���5U��<j�J���6�<Z���v�͕r�v��s��>5���V�ނ7GV���$Y��>�:�$z?���o��7SjY�y+�y��wQd >����A��B�k�ҝ��Y�,7~���{d=�K�R��ɔ���D�Ғ�:*(z�ߝ��.w��|��&�a��T���?�a�v~��ڰs�Y�Q 8���TZ���q��/����3x��3Mռx=|ڼ#\��9A�v�����[H�.<w����k�}��&�I���G�ZB�8)�������B):��I�������h��� �=���f���`Ñ!k�z��9S��S�5�b���֑̿8�������J3�e��	{s����|��<:�u\s�p����bE���P?Vzƀ�g&����a�X��4oRa�ak�2|eKd�VC��:#Ǟ�l���+?�Zas�")�ma�"�sN�0�.8?y��<�c��ܹ������/M��������9�k>�P�5888��i�}М����X�>�F=A���W�e[�D���6x^�����蚶��{�
�1���:M:8�]�h8bN�z�+��q�F�S���.۵�6L2�Q�[�H5F�3����̐o�*z�o�������c���;�_𘺿촎̬lޖz�å�6�{R���Q��@�����_�~�Kҕ��[�7���0�Y��z-$�5���ޱvt�4��%g׀� �֫Vמ��@�(�1a��y������S�J3q�I�Ԣ��j���O�#�����2048���B)���$9�o�u��f��:;��|[�'&�n��Wg ��P�yB�{g��� ���6`�$�#\CZ�<�>��v������a��v9ׅ����T���a�MZ'>c!ݵen�ǝ�.L�t�3���F��ɉ���EՓ��`J8�7������KwV>v��Ɇ����7��8�"�r0+#��_�?u<�`��eõ*W3�.:�h�T�/�d{_�y�Ŏ�����@��OhSZ���h�Cy���8�`�|m��T"
�I�_3Wi$�So�_�Z! ��	 ��5n^��=��A'dW�@IӮ�c�U�L�]*�*�Bl��Y��[%�K:2��b�<X������
R�b/$��9U�y�xL���c��9�)��N�ꋃꉈb�	���Y�P�ߚ��*�
]�{H�����s��$m���#DY̳i�~�#�;�SG\��ܙ���$�����`�ܒ�'�x�0���Ir�:�e|__��w|��<("��{$��k^����T�}!�MpV՟�st�#��|Km8z�Y�iP'N|X��~��;*�)LM�N#�hf�p����7rp\r� v6q��x��O��X����������_��J�U]��q��jʕ���%�ūq4���B��V���`��9�D���l���#(���%�8s��b�����׺��:64V|��s/Xe�N�|����|�8˄���:�ݷ�U�WP�[���� �='a�ɥ�ӇP��?w�A�d?P���µ��<%x-�{�i��Xdl�츦V�b�q�'����<Ԝ}��?���N'��ʤ*��|iq�K��dd/oB�������P����pE	!�~�]2�/��"��S-�z� =�ep�R���L�mT#[��l���)c�%�GH�ۂ1��,I��tI�Ps�Ɩ)�K�n�++���IR������+|2e����w���c�)�<����f�t>�Rb��NbSy�Ş��0@L�y�9h�L��I�-'d�������6��ۜe�co�;��"!�W P�2v(_�V��lma�����b���$�D�~�B`�+#W0�ҟ��Y��B�i(A��_��w��`F���*�LmЭ���H�-4�@�QT�����F��h� 틀E����^��%hn�l����R]�t��j0�l�����Q-QC�WO�����x�)��ʈ���O=�~��w�;��wF�}�����g��Z|~�U��!�7N��c��<eI������W4�[�%`p!򫠸���e"��A�/g�J�xV&Ѿ;�Ii]������� ���Ǫ�f
�!>�s�W��9y�䮸�M��e�j���ע��]�*�U�P�&�¡��A�\`�x�����p� � �MK�� ���n��VxD�g�v��2_�Hh։F��B���]��Kכ��_Y��z�����;{M�"/O o'A��	h��f�[=��$j��_�Y���9��7_���tD����%G�C�l�iA����Ơܦ��Y�W��t�jL����L��r$���Q�g�0��|�4���D5@4eƏ�p�0q���cZ�� ����F��(����m��>m�{gB���"�?( :�7(����5��&�@�ݠ6r��f����ד�id��W��k�T�^9%���p,�6�Ŧ� � 4[!`a���4�[�����y�A?�d���l@(�˳�������^�}^�<K��h�i������$�i��r��u$d�|�|����-��ؾ�V qr^�dea�j,�V��lW@������ϻ��͊
\�C}N����^_����{?n(��k��yW2�g.!�A�?	��l��U�'�}�����F��E�[N I��)ǯڀnG����q����8x�kv�t�p&D�ӠK[��κШ9�9M*�ϙF�b�	��i*���&��&����k���Z���l�ӂhm��q�1�}p��|�Y��EsVK������r^��`?A��y�!m������|�}��l�5l݀ӂ^�C���:+�@AU�d�UŇ,�VJ'Ɋ�
��4	��*���4��}CiXC�/�r�!��G\�t���e�7�@"x���L�U+?-��0}�L����7zBZ���4A4��N�L�2�̇[�k��5BHUG�=�#ߴ�xJv�-qh���UH^���VQ���ms\��3?���;�S��iWoZ���.u���U�?�2f`ۉ8�U{����9�I���A����ߪ��({uYu�@������eFr� ��i�٥�T����ѫ:�:�7�3�j܄ފ�%*s3�,�[�8m���!@�s�|���>��y��9�=;RU�����a
�|���8�ۛ���2��?�$�OK.[�C��d{1�^��|���T��z<dJ	��H�.��8XW](s����f�S)��R��ot2'�i����"��-���g�jxhTߚiP��$��V�5i�aR������F� Wx�srVb�q��k@{�1�����z�A����sׄqx�a�R�������TGlk\NZ�Bt����|<�ɠp��2@�g���5(��f͙,ݴ�0��lPā�a�?�T���d7(���v��S�\0V�i�j�F$~u>Ow)���׎���*�c�V�c�@>�"]x�����fW�<��=u�@J�����ح3�t B�F�!�����$�p����~��l����g�w氢�85ŋ�����BLG6G�U��&j4u׹>���=�a�(B�j���I�F�Z�[�t�\u��_IW8�
����L�+"�Aān4�S�m����ne����վ��UO7�֘�u�;1s�����|�ҭ���hw������I[�W�nB�QPS+%�֖�t��T�@˪cE�i]���D���ѡ�N2Q�C�oG�8^��.��>����l��W0@>�O�_�����ǅ����Ҙ�#~!�dF(�1���h>��C+��9�����C��2Q
@HOA-��[�O�vK=49r��Ew���m)�MɊvk܎�!ј�m�N����a���g��]Z�i.��T�r ��A����ͻ'+|��'`(�v�X1�}m��nh��[������\ӎ���W];
����_�S��Ќ���|������->2���sbHȶ�k����h�U�}�r������U��랚4+�틷��Gnm���y3���p�������U�!.G�$��޵>�V��2�
����/1<�[{@�V�f�}����U+U�#����O\"G�%���Q�.�M�f�4��rМl�x����tN�M�tga��0�j�RĔw%J���[� �������Z�t��h��SGGm:8݅oJ�zY-����w|����e2�UT��� B����Տ��\L5}FU (N��vc$�?N��W�ڭ��PbFK?�+��f���Wש�"�jj��ian���~
����N�N��MZg۩���ͽ����ѹZ`J���ol�&��O����c����CK-������l�����Eq��XO�,��1��呚\ �JJ�o����޲f�yx��(5�&�2�;�P����!��o�ﬆ�a&��^�J�f�"/�-��cԀ�I�5�+2�f�"�?kK�z�&�N����JZ��05�|�U�����e��)���"��F#V�:�50����'K�I�s�V������t����1�&�]?\�[S�":=�4^��3�R+�\I�5���L�ܲ��&W/�&�"e��@�'�2 ۢާ$�|�0LD�Xc�Q�wYB7����e��BG�vo}(�Yb{�~��Z��#%�b��[��������q��&h+p� M��@����`���E���ru�"O �2��m�F��5�_�-W�;���:INo�@�I��$�09jז�鷗�jYj��s&]���*��
!�xꌰןS]�S�>r~���r&KVx=��X�|V���ݡy�BV��]��� zT�0�W�YnR�V���U�Y��U�v�N�B�v0d��L�II�on���eh-����fF �޻S����dս':�?���{��Pܨ{hb� �mg*��q�G�;˲ŉ��y;��,�� ��s#W�u�=�3�V�7&���w��~8�m�I�i�"�	m#��?2 `�	��2���p���Y�5�~�ݿ��q"�9����VSk�!���hjo��>&~GՌ�	T�cOmf�n,Oa�1�����<=�,��4�S����;U���Wc���g��9��p
.�<�?�^&�V%C]Z�ݕx#v���j�84�bƸ��wGiY����5~�������#�౎N�O�ƖE�ּDnu���|��:l��G��tv�K�����m�S1��>]8!WH�ġ	�⫽^�7޸���|Ct��I1��"����H�����"'�pv�6��G���֣�)r�P���A�_�oe�36ݐb8�����Xm�=N��éI'��jo���Y�nS2���[ۄ����[ӷd5�c2��}Ϛ�oV�C0R�m��\�i��܋��f������a��Rs	N��լT�)��g��3��m'$��!]�6.�;��]�2 ��v�u�iE@&J��N�v��ǲ��A���ϰ�I
E@�fW{�Ö�=��V��p*���u -�i�y\#o��-0穢�k!�ns��2��.9�5�K$�d\���K�_jtnj1ev�S�T��b�_$��+Yz���L��i~���ֈ�~�P���뾅��fXT|�Ͽ���$y`V���4�f��!��쟲)�O�Su���$�=�ۮ��(q�����$��(L{��Lv���Y�)�9�_"� ���?�
�
��N<�/�}lZ4��(DH�ɋ���&9Si��]��"��/��`�%R3��F��NQ���g�2K�!���E��#�/6�|�>^����M�2��8�����G1�v죎'�,8����37dV�ʡZ���]ܥ_�{|��ӜU�s&��fV��������T��P:�L�v�M˥K.Vwr�+�?�����p�6�p��a>� v���RxC��;����}��30�9鰃2x%|$u	^��<�ǹ�k!��K�
��@�˸�6.�{�hq چ����Z�?i��#��սKL�E�����]j�Ñ_Y=3Ir���_��iu�9�3E��|~��w��r���˚�x49��n�*�"�x*sx���CL�HY˩_J�@���5}_�Z�ی 	I�u����n�	��t"�d~_rHCz����U䫋���4K��I�S� ���Z^-��1��-O��*'�lu<j�©߀�4�bY�	�D�%��<5��v��o��d�����IaaQ��k�7+'��}x�滪m�i�B�gU��X�V���#��"��4]�'���]����-l��n����w�#��>Y��L����z����_�U�Y��ԨYT��� ,�s}�U�P��w�P��p6��s���P��MrO��4"�r)�ѭ���*��dـ#��$���?�	+f {�A,�俪��A�;�`���|��u�߸��@��߹�E0��m�=�H���+�	)��1�R	J�ŕ����g���Ց��4sJ��v)!����B�gAR�k�+�L��S�H�d������q9�����"*��Og�Mq���D��Z���e�B�l�IrP#�D��a��g&����d��K@�'������h���A1�.Dd��A���2�h�1ً&����̞=:A=�I��f��Y]��9_Ԓ�ӑ���W���--q��Z���Lj�^Jw���' ���:��:����W.�O��@=������.:�=p�ڧ��Ŀ��ENN�T� ��u�=��nc�BV��[������� A���Ud^�H}����Џ$�#)�wO�,qZ_�I�l�_i�=���M:������/F[&X��I��V0���,TY�W�?՞��p�~	��G��ˁ�m5.ytGmK_�j՘�x����A^���|��t�����@h�k��r��/.B=�p/�ol3�YZ����%,�[B�#�K_�F�����7�2���7��}����2�7`��	�!�Y3$���?���h���/���Y��.� jb��tG:wҷ�^�ѳX��Q��b5iX�A�)���)۰����4JD� n���@/T7�n`�	���=�{N��@tX����8���hv�-D��3������;xZwŁ��뼨1��9�i(�܄^Z�ed1V~x��f��(��cfI�@C�h�Mݟ\�͋<<�X��SUѓG�d1l�E�3�O�	LT7�=l�����K�I[����,����f�۟�:�����}`)�z+;�i���퉡Nf���&�G;�}M�{t�_�����A	*qv�Y�_��S} �7*SI����^�_�!���8Y���|01#ť��Gx:�z2��o����$;��;����Q��kRl�o��Ei�tg��;�Mq_ ��g��d_Ɓ�ر�� K!�f��� �U��io*�KU~W�C8~إ�?U+ ���B��rܷ�Z��D�I� [ر#iogb��((��9�̄g�T��Q�Bm玐G�|F�>�'fm�/9YQ��e��θ! ��#ЯԸ $�ֆ���ʥ:�O'��ӡ,1�/��ß�2�c��r3z�g��C]��%挩�b�)�ټ-�r��* ������"��>����^�TZ;����:#E"fI���.�w���c�N������,�̇���1dM

 ��xT�>0�b$�����=�$�+q6W�@\ֲ��wk{_�,��pn��?�/�1 ���Zu+NG���\��[��"p$%�B��(�/r��A�;(?���U<�?�)	���AĔ�E���0���T$��P�혰qJ��K�dkTZZ͒��$+i�t�aU5�u�W�ڒ~�8-P��8��Fh��G	��	I�����1���_�x`V�=3��2��`��w��C�%���J:�����'���.��p�{4�0g�(%�>=5/$��y+���kW%�&��,��>H�W��[�!�V�ҰUX��������2��n�qї��?��{�o������S�Ɓ>d�.���c��N�C?D=�Sv�!_�dh�����|l+#9�l�#+Ge-��K̈&mu���iy�!�|&�ܛ�n4"4.٠����)<`��͎�PZ��+`����������i����S ��i��1_�;�uKЏ�)�t�����!�Y,"S,GE��+��n7���W�T$�	!��3/� SWU�R�����ك�-�Q�k$�C��$saA;L��r�ʬ>��%x�Q���1�2V��q�'OM����+���&��G�ƇE���#Ǒ[ou�oU�s]��ص����\�Mդ#���GC��&���G��)4���A�����g�.��c�����J��S�8拁��])G���^u-�l�5w+Pr۪c�2�#{y��X���pP��T���G�evX�Sܿ+y�Br�*CߦM�>w�n�5�Efp��LR�-75�O^��ʫ�T�
f�s���q M����'���co��j�Ϭ=�����'6�eI�MW�a��G�|�bQ�r�YD��d⨀э.}�@�Z� �(X�@9q�� :a�{��@�e.Hx�cl3�O=o���po�:Z4l5���Y�?Ϥܶ>��[-p��I/�6�߭��£V��M3IN���6-7��3�u��i�i��� t}N�2���cB�Щ H���.���m`s4�z� ̜B�N7��V�Uŭ�5�NU��F�ث"u+\"N8B|�u��1������6����!Y,B��	����� g�ax�|�����P���L6����fw��@�A�mx?� �(�.{]�2�jM��=4{钦��t�Ϧ�#���j�=�Ѓ΍��Z���	�������MM]����x�Â�&��%v����Y���ތ�A��Wd��ԼhD��.0D�63RoW{�î��\T&�H��Wʰu�d3+��;�Qö���|5d���B�Z�5�n5s66*9���u.4�����t,��1V=��q��F����V�������-�1G�������)�c	T-@⭘Piz�d�hA v�G��'���CEgoA�!Hj�*۸`Y�`�N��~O]נ[c�N�D��5 ��	yܯMy��j��g-#}�,K�!OX�m(7xPm|&�ҿ~�b]��I�δ~mp��gf�tepu��v��e/�@���]\f٧�r�|�m�?�uRu��<_���΋��A}��"T��9��V�S����.Q��{�Z�Y�ݔr���<�ݞt����째o����2t���EtI��x���>��x��َw�ғK�~ ;�AM� ���E��[��0|��V�&CeM!�?e[)?j����f]����a��hDU�����,�:WO����T��M!5�.v�J���@qKIv�Ep��T��H"ְ`y�j���8����������ǂ^��b=�x�������ǔ&���^���t�ܮT�4M��3=a�J���In0��I=�����Ν=�͋~���WiNM5�8J�x�1{�yl�-x;��^ċ4)(��0�ȕtUWs��D�[�[9)(��M���k�g9U�OY���,��bf�״���S���ՉJAhf\��#�ù�B���2,
���~F�z7�U ��LIyE�*�>����T���OqP��Z�=45��٣  �D_�VټE� )���[�Z/�1�x�$��`��OV�S��A����K��<�ҴF��ޢ](�!�Yw�߶�m��Gv�q[~{iuؾ�u�j�����ә�$	�4�[�~i�L�(R�o*��)�:2�.)W��X�s���ʲ�XԚ�A�ţ����iU-���zA��j2@���N}�]B}�4����V�=����Zm;O��sP��+L�>}��N�O�y�����ǻ[��y�a���6@֞A�˫�wLh6e:",T�E��_����ܝ/�U�},�~z��ʦ?�h�⣢U�85��PW`�����<��h"x5�uq�b7��zO��a�f��wY.��G��n^��|0A_�A^��Z���ʅTq*C�En����YG� ����@�sߑ�r��7��9I��d�3�t�4Ä�0�ݥI�A-n�c�����&EP|ʃ&{�?� ��, /�Lr%,g4����1��1j`1�8,�|���󩜾]4����Im�Ҕ'�����-�<^�'-w��ī�m���Ȗy#h��Pl��N���+���.���>s��}�2�O=g~"��hz�[dQ3�������e��x��Z̿w������\��.��h���mR��1j������ӝ�F�J�/���]��-�T�"�{=�"-!"ȓ\����M�a{ȒO����@���o��o��`^Ggl}+���.�Lp��d����"h�SXq�.�UD���Ì6YgЏaĨ)CП��0=T���;�XK���0��ZT=Qfwi�y0L�ѦkK��/J�i�nٹ�^���)�6�{�b�H;Q�A?hO)��@Lx~���,��X��f���W��=�s��JAN�f���5a��8R�g+�-��޽ �����o6����xx�X�bHN��L-}���ڟ3�5,�(�3~4�8_��铋�Ri��?;�Q���#y�Q$�+�����ݏLO��y�j"q)�?�E��u��!b���^
7�0�&��Ko'��O&@�������s�z��p���.�u�~hk�7�x*IČ{���(���k��+�$�+�l��c�(�ےx��{���9K��ѳ_���3(�E����J!��J-#.���Łl��1�WU���v�L�/��K�,�����`�Z�?x�q���J�tװ&�;K��:̙��$�GU�f{<s����\Gw����W^��Cޜ��)?hEx����h=p��<���w���gӡ���g}͊�V_�q�SV$���sU�2��ځ]�>��������
���cq���W�0�ɢ���?r��$�d)o�,g�2�^�\������I�ek}�p5�<�$���X��7W�bV[��⯋�*Z](���fJ��`�v.@u�I'ó����&=���C��5�
�YܐXAv�<�7{NrC��(.��U�>��f�Ճ��"�c���\��ƉYuj�;�U`���fɤ�A�
�����l��f�V`ʡjw���Mٗ�W��L5f�� ���Y[��z�r�MA�o�`�e�)ω�@����fN)��4�R���=_����w7�.9zo3�t��x6n�A&�o�1qW�����9��i�Qʍ�0�s�d�p!�5 r��)E�ti��tww܋yq��_���P)�l'4���AJ�g�g�+C�'u��&��h������7W�%!�x!I����-mYF����YҺe�M�C5v�#�w9_
BE�^����J��M����4"e�2��G��{�����@d��
N���- ��Q�o�}p#�Z��x�F�Wې�4�����B�&�a,�=0�|�ըo$��7�H��ͣ͟��^3���<�7T��x����l�qj�/�`�e��>g� �F�r0�l��)�C]��Dp����Py]�Y4v��-f��S�/�.� �)u����}��t� �nO��c���׾�P��+�]W "w���F��,�*XT�SK���^���Z�1�t�#��:;^�T�_���7?�7��S֎<~���*)�(ӊ�V�廬�#��-Ěo��j�{X�_?;@�����]:6�5��C��5r,>PB��q��Y�/Fn�p�}������=�-Ǣ}�&�|��_P�]�~����d�Y� �1�!��R��g�T|��-�o]*�Z4�$	å�vA���P3�o��ѵ]z��T,�z��!�x~v�=�q쀡�D�wv�I�x�u�wU���s��@�߇�Sۉn�[��I5_��e����I����֩I�B�Ռ�"1�{��i�=��3��}
�2�9;�"R��u���*�}�����J���G"G.LP�vR����h,4]���]����h:QU��B���h���#)׹��MߋO����<j�b {'ǭ�zG��#_��O��A��x����a+y�L�?���<�Rp{aT�V�J�

'��-5�G�jY�F��sBbwϞ�C�]�K=[4�2���j-���|�Q��P�h0Āq�F�}�/�
>}�I���X����	�+�a��8�wd��W�4�����q�~A�|;n��d�Q���gc΃?��~���౔#�D�H�i�ye���~Pߗ�[��XUi���hT#5��8!�/�E��("\�������6BK`�:mLpۍ��E�����3F��S@�3e���/{��ـne�.H�D��X������aj���=Њ�O�#�� ��\qE��%�J��\Êq�ďj>����I�-.\�1�S<Ѹ�a"|��YZb��e%���u�,ʥ�Hz�F�ԩ�E�2��:P��e���Ń�M�5��NYtI�y(~�t睁�+M1���=P͵�Ϩ��r�Si�ro��`)��Fc�k݂������eF�X���u�&c;~�Y��o+�ɕ��jj`%�oK �)8�+M�h3��sQ�0��QT9K��+ғ�7�������)<�K���pQ3	jN��X��쨴�Ł^������v���������u[����b�2���#UP"�<�s$��[��5��\-b; ���`��]��!�h�q嚾嬢s��x�C�Ņ�L)�Qs"�<Ț	��#D���{�:&�����R">Ym0r�F/��@�B<{b��fs-���N%�U���:��W��,����+P0�&�-��ܣ^i�%��o��$%(/�������q�����!%7�Z80uX�e�tڊ�wgR�<��U)<
_´����f��+�\BvU��>k�ɭ$x���%(�ܴ��:d���s�!\.eH�?d�TT��<������J���)��ݝ"5tJJ�p�ni�nɡS��������X׻֜���o<��g3�_�|�҂-�y�Q^	��.LD�l&4�e�pf��i�{?m(^9Z�(m޼��w����-�	3yx�����^E�I�K6)Vq9X��S��u�͉Ŋ��wa� D�~�r�y�R���t.�<9�m�7̘�0*�+�k�v1@W����W=�d�:�
:����4�o����M4�P]��)B�B+В�_�2g��n��>�w�<7A�ڱ�riN��$2�N1����f4�ע���bA���^��o��2A�Ľ�Ѷ��ܱVɳ�`��X?ê7�j�/�����${�� -A�'�� ;:m��=8�p�0����%w���8�Yj%�Y�|G��FgDRn��wN�+�o�a�oO7sLg�ژ���'u���� DZ�������2~)��O ݜ�Iz%X3ZH�iF���q���Cw�\�����p+I�������~�rvR1���RY�ݪ�$[!�i��t��o�~�ikQn=ڹ�M�7��H���&��짹݃�=!��ǚ��3��y��p���,�n�M��HZ�{ʺ�����6T���m���8u< ��+�7ʯ^ŲlL�P4x�W����M̎�|>'d+m8v�$�-�X�Ryp�Nb,K��s"3������D~�ޯ3��߆�J@cִ�.G߷�e��R���ؽ���\s���kw@�)z{Q���N��R)}F��$E���j��axN駷�C�h&��Zj!ʒn��іձ�O�&2�d��<�k了��SMh�P0⤆"l�o��ZOD���)�U/�s�G����׃�F��/)�p��-E1N���9hDؾw���n���E�h�	U�\nt�U[Y�I6����[שKf�U��I_�M%c��t��F"J(Vu���fM����*�dB�����
s#�m�v&A5��G���e	���C������7�k�M�.;V�ھU����FN��A��a�_�x�eZ��hKa.��M� ��w�p����:��i�j��*貗=���J�ex��̅tr����k��o�^?5��Y<q��R!�(?.F�!�u��j�����Ȗ	̙��=ƍΘ�Oϔ�X��zG(��oD0�+9��6[�%������v,=��_�␜�|?n{:]�4�锭���ʡ�w�; V.1N�ǚG䵖��G9Y�_��/�aj��0c�t�1�?Q�Ի��N}����xF�P�|�9Ŕ7)����g1u.m�o�)z��:���yUC�������6A
d�C�H�׶�:,�~9����M�>B�H>vp�k̒������;¡�ܱ�|Ĳ��3j�,YGX����m���C���.ö���ύ+�^԰��g;�<!^�u��/PC��Q(�4�hd��{+�q�K�9�z#u��C(FP��W��>�Iy3�,���5�$�s�C�8�D�J��*3�Iݔ,�����Ϊߥ�gOx�L��l�O*pd%�_Gƌ�e]4�d�N�vZƪgM��8^^>��3۞`�/�c���
�^ŖS+MFK�p��$�Ձ�W�r��"��*��K�Ŝ��4_ΘU�+I��D'A��We���Y�*®VVB�Փ�[I�mo��c&?�A]Da���n@�v��� E2qm-��Ky�����$���&YP�SaRD�4J��A4�s���ۮn&fZK�\r��|ց�n����ec�����n?�{�/�7WQcz|5�!\���ߝ����J����)���w�֖`C&�R����^stD�O�'�q����~t��ć�P4�K�?Н Ꝭ�5��jc�$F��s�j�Nedf$ϭP���c谆��g�|�[;.ME��.߹߄' �;�C�����X��h|dv���x�=�fZ�P�6w���[}|��#ӄ�����p��P���pO�q�Y5ϭ��^Awǖ��p��$��^V��#ޯ���xQ��ǝ�u�|P*i���َ�4�����q�'z7^z��A�(W���e��	��㎰#�w��ku~`K�`6q�'�5�[j�p�����Q���"�����b�"�׉�zᥧ�f�r2�>�v7�f�C9�ii����ry�Iz���e���3�Jn���:G��
�K�S`0�N�I-��`F��K��s�J�V���n�K65CȤ��M���Dje7����������2be�+C�""yh���1������b5pm%�B���%�j�����	��-}BK��j5��'��<�����h/�lq�7�'D<�7�kb��S��ll$�E+뇭����Fc�a�`�Ib~t�t����oU�����Ҙ�A�,IY��uSjE[_j��c��x��a��.�kH���D���yԉ�;��Xэl�H�Yԗ�<���JV~J*�(��z��A�O��=x�	�Տ�e4?$m�Q��L3�Ji�Q#1�g����?UUH��D���ެ��sڭz�ͳ{�˗��:z?�<N[�E�u6��[��iC�H��.Nu ��đ�«�ବ�����=c{X?p -�S�b��ZD}�^!�����4�)&��b�Ɵ�&�+T�����d�j$X��Mf*8��"�M���v��S;[	\�ξ|^��Q'PTEOSc}�<J8%���y�� �ZW~���;�ιn�xI�ZE�k_�n�y�h��$_i�B��5�%m8��P��(Vq>�+;�-��O!��[�{��&=E޻��7i�d̿h ����h�����8Mrz�PC4���=:��/�����ď����:���<����sŇ��3�\J��Z+�;-�c���Ƀ{0���v�P��6�\~���"�\ٷ���(�������˴���	O3������2�����.	5 �nr��l���C������'1��\�{(����&�M��E\��^�á�l�����-X��8@:�~b�{��N���zb:��(:�pGE��&W$+�Q%���nHW#�z7�Ԩ�C�F�tE�΅�wO"�l��ն�mA2��zY	�i*��	)q���R�����>�Q�BN��`�a�vs�40�c��-�D�|V�+�D�%��Қ5I4jL>)�[K$:x@EvH�u��skl���V������G�r{�iGG�����PQ9��lph������v+HTs[8棆[i�;/ܰore4�Z��#���[c�/(%j��,��Dz�#�Z^#2��$\q�Z�!IHJ4�g����b�9y�e�it�Q���!r϶,�u��gT��z 6a.�X8���&#��*?�a�-3��eCZ�o�����1ޫ��D�+����ߠ[��a�d�G�0ȫ]������I=��#~{�4ls�A��R|�q$L|U�q*-�x�oU�w3��Q��P����G��2���K&AKB���3��;�_��xv�^��-����z�Z����H�nI0*���syn����@v�p�����~��R⦒���仢Zjڻ�?V�x���va����s�����N�&���G�<��N��ToH���2�t���l��t�J�S�|�a�c�Zio���0^G�{�H�
�d����udk�R�������K��J(�[�^�:�zu�������<�g粆H��ﱵ��`O��g�$`0�}I��ީ��ꤚ�ُ%�q�����M�Q���Si��K��U��������+a�2��0��2�R�0Λ<�,'��2��\�<%�C�;�1�'�������̀-�7�ϙ�B��;Ff_asԹE-�>�>���7U������G��l4��:C gUU
8��NN5�<펜��$6d�WL&��Q�]�����r����Ar��������B��(��+���5U�gf�H���$�r�uy�@��[n �	������jP�]qws<��6q}�[3�hg#cz՟�55�iq�t����_�r���X�l���"j2zyB(�5�o�$sr@�����t�"�c���G%�-Yp5�\��v�}���5=�6EH�A{o�Z��<5�Yp��,� n��3*,�M��W̎.#u�S7J�����:}%V#+�'D�֜�2c��:$�*V~��_�l0�P�L�Q��j�%z�g@?Wi�.���� �Ϲ�`ܑs�:�.S��!S�G�I�|\4�Z�J�$�xYl���0C�6W���f=�	_�B5��&2�?���	��E��I���^L
�E▀�a2�Oz�U7>�c�|.�@�iV�r5B_c^"�.�4��GG��7Ia���3�^�൦��*���h��h?hJ��|P�x���(�D��Tf��c*�P�ɨf>����8��u�<<�ޙ}xFM��������&�e�&���RF��=���E謢�ZR+q۾����V�����{!&*fD�_�qp�������7��UF�r5��݅4iǸ�

����|J���?�J>�cm>�z4���n����	�����%�I2���a�t����y�b��8��c�fCE�XH�β9ޕW��!�^C���t��qT+��`^��[Z�b��,G��դxΨhzӕڷw-'�i��H`���v����AΤoR��{ϧ��f����.�TE-G�������Ka>!o;932N�-��,4��솫�$�����|�c����I˰����\x�������y��M��r��a���)g�(Naa]ZK)ZR5�}�L��<	�Wr���2�g�^:Z�qX2=�F3�b�t��r{s4�Z�w�H�ϳ��4�tRF��5_jl]ײ�׀����l��p��F���ˊ6�yCέe���RK��7��r���1|6��	N_:?�,��@PoTg0����QA_i�`��Xk�,󈓼G>ږ�N��A�},�n�������LƮ�����L�t�����f�����V�7�>c�D�������i��i��r9����7�d_�{���A�W%�Yu�����/��?�ۅ�vv��9�� �Z0�r�B>{���w��πV��`E��(p.5�x�N=(�s����*?{8PP�O@�)�df��W8����*
��y����0*:�}"�5oS�/ �ӥ[�퍍�#�穜���߳ 6/��ku$�`���]�r��Q*���	K64�7����Y���g�-��͏]��7o������9�Կ�FG��\�E����x����*�f�/R���S�04�n�cU�y��n�>���>6�Յ���6��-�('0��󕭺��ʵ��m;������0
���\�mU�Pj@(����w�Z%V2��0��bq�+�;�+�{'{9Q���s��iFK=�g�`�}��Y�E�+�[{I4��2R����a�������;��&��;4� �n�c�|W��eN�hf1V��X�6�E@����zC^��bW�Geo��`���!0U��zM��/r��e"���l>z$�%���%�ݶ ���o<ج2�?�幡v��׫���p^`���%I>��t2��)�r=�����;XƵ17o�Z\ܘ�!D��lR���`�?���RSe�x|X�I�W:�@�(}e֎�rT�ww�5��@X�Ɯp� ���z|Dڕ��n��
���i�����hL\	ZKY97�M��QF�F�M�d��=����*�>��7�^~-}�.k�hcf�P�]]�í��P�.���҇��Q���'�)ӊ$�9�,忞ֻ�!"vh�g�v��@cx�^�O�@��h����������S�e����À�Z�7S�&���_��aԛ(��M���AcrR�{/�$K_����);N�Y���HͭS�oI`B�*:�e������ }\�o������Ǯ}�Y��V�=;7���UU�W�'.��h��Ӿ�N7�B�s~��.x@�:A@��`��u@8�/S�������E���b������H=c_�͇7�� X� Ǐ���bJ�	q$�Ʌ���=++�:��3����3�����;w�~����ËOH�ݱlkHI�������Kg�lae�侘��l�Xx^�k�1�Q��缴�e�,��vF�-TcGk���j:�΢���
�<:Ȩn�Z2�c��ږX�>��%/I�KBN^�����D�:���K�I'`�))�͂�Ϟ����b��fbeU���
����j�]��6<�����NN�ii/��׫���Cz��7OyE>U����y����D�:::��f�3��`�$��M�m�d�����ۑ�bY�C����,k+id.)l�����-�㓈�@<�� ���-*_Ô�5σ8=;n����
�G���/���듐���7�����ə��Wcs������] Ԋ�:�Mc�gihh����l��h��x�$��;���QM"/aZZ1l"�/>D3�͐��MIi�S�Ml5W���/%��v%y���p2I0J�W��^�o���?u�Q+�Ac����J�M��k�]w����lnFƫ,�dU)��ɩ)NAAK�Q����j����.If�je�pc33��s�R��$j�+�����R
4+���'&r�CP3�s*RR��1�L݊t��ņݥvK�ڞ�#����F�T9�4Ji�z	��^
 ?�| ��/�cC����RaU��l��mGӓ�!S��/�M�Iʒ��ʢ��n�{�����\�S��4��-��`��{�!(_t!���S5P\�_�8�����;I���dRf$��fH���h�IfR�u��br��~����n����ְgܰ���h"hr���� _l�v����$�<h��v�<O�$@&j��E�h������&n{��ϔ0���===|��8B	�!�q�::�2�ܜ��w�f.�:�:I��Zu�+���/���ME��(W�Cs����~�1�o:Nj%oe�\�+��������1q�+*�J����\3��v�܎UC�87�i=-&�u'�j�n���i�~/?��N
ΟI�v�E
 ��x��.z|�8�C����KI9�3�I��X:��TG����1�U`j�?i������|�\�D8¬�mZ&���l~uy-~zz*ݾ�Q�aJ[���t���h~Xr��8�� b�__~���u���l������Ǵ��f�M�U���d��[X������,=3���NQ���	�N�`D1
�S�@���C�b�Ľ�}���o�bd�_���AN�t�n�''ff�XN��f��;Ϻ�͝�K�w��o�~n���luؙ�9]�"+Ӿ��Ťy�H���TnXPq_iN�a���l�O,��62��E�In�%<<���7�LF���+��d�%�c��l��W�&�y_y����!"lIHH�d�M[>��pkϿ��AYb�KCCS�~l�9^􂒒2s��$�j�����(�/���=��|�˟�@�iE��#�B��������M����t��=��1�,�@"���E`<�J��`m8/F�vY��102WLմ�S����\l�0�uf�yu6���S����#���2��i�L��:
Uf�Mh9[�Efċ8g.���$��騥�-�*Xx���yG/���[�R^�����`ʏo�&1�q�yo=JMG ��z���9�D��V����QM뵢vr���#6)��⨢a$��߸J(h��r^���6<�yG����*��l�d�hvg-����#Ҕ��<�=Bjz���q�=��=z)�>�?nx77?����ۢ��d�k���r�Y���KmEgܷ�r�H.8&�4�����[�����o�ؑu�8(��:��TXN9��B�x�{Ks�h3�drXZ��	��� >P��oW�u3�fK2�Ks��R'#��"D8�Gt	L���>�B��!۝GL݃�cZig��***����B��5���l�`c�:wyT���%��`��lk��]�J�[�B�}��S��vo��%���V�"B�:V?�蛔T�^Q�^حDe;�0���A�؅�T#���
W��u<==3��~y�شܭ>�uWQT|ˇ3��o��%�5���u�m��=�^i�T�Ed��W�'}�:�wp�1`���So��9ha��ݩ� I5��r澸��&��9h`�P�ȭ&`,�k�12:��A�S:0:������̜�6��syy��{x�@�W�N���Cݫ���m�X��������^���A̐3ϣ�du��5��m��i}����
G����}}cDb}�&�1��:x�����+�@a&�Z�?�w���.{wE4<x0 �I���V��-:f摋�B�ºh�9�p=.v��9�&�����LA���
��z��x����]Ջ��[�x����J�44�+��~}<ȼ�zΐ������4�Tߍ'�����g�g`j(�����=ܤ½m9W��Z����@��x�Rw�[��3�}��]��&��S���s7��ح\�}ڞ�j�_����!�|q��b���ҫ9B_��ئ�M���\�x��f��?�U�L��w�Z�Ԕ��v���䔗�VUUe.�5�����>U*++�C���	�c;�yU)��AhN�b§ak����.�Jc���,��:dĞ��0k��^�m�d��ܣ�\oz����asޖ�GLf�8�yhѶ��to9��O�Σ�����חA��n��8�v	��z�	��5dmN-�$ԅ3Jx������̴F����nؾ�U�rP3w�puU���=�R+5�ą\�U��/�3�n)�t|&�nW��8�?(�`7��r��O��8ņ^�ϟt:�����F����r23Eyyy3)o4����[N��Y�a���R�y��O�bM�dJ�{c�AW�r7D�ou�;:;�څ/� �0o(o�u͂�н��3�dL8�!u�n�B����vǑ8y�v�"�ܼ��o��;J4%%~��}� INu���	;�$1l��"�d�g��J�1l^~�BMS3���0Pcn8}�����OZ������H����$Wѡ�!��4J�u/���چ|X0�(~��ZN��3��'ȴFC���&�_Ǵ��lOSÈ�f_�� 9L%|t�x�$�	���Ղ�q~�2` XXX��7}����y���5速&��HŌ���1���/.6�8�ac��Bh&(��_�,� �,-�(Z'۹��n�/tҞ��Z�$�,:"ęs�C_&#��O����V��t����b�zI722r�s_�򅤎�No��k���p��r;�%+�UO<�ۯ����-�35jS����*ۣu��q}b�'pr��ך0)��}6��t�䜿{��%V^�Ac����C�[DZ�}��ncrb�["�h{j_j_K��Z��ly�%��À ���J�ڑ�5���u�~Aܸ���咮���W�iz�W��s?^��M�g"d�ٯ@�g-L�|���Z"V�a����M�A���{[��ksMe��d��2�DVI��j_Ey��f��n��;~�~���>y����l��QF]qxe̡��剜�BX��������-***��6�]f�v�bSX��<o�n����!ወ�_���H���1��nq�A%��f	C����LWzA�IJJtP�d��69���I�~�{�yv�I~}����QS<%�&��c�U��ʯ)���7r��(=�o�T8�E1}�����a=+i2[���Ȩ��p�� C)KvM��P���ˈK��;��tzE�]i�Q_����n;T��i>T@*7\y&�9v9໌��f��[��]n�A\*X�&����f)BF��A		R~�o�B�m�$[��po�����P|�K��>B������6��T���E)t�~7f$�a��"��А��^A�v��}]ee�6
f3�$�~�O�.L<�����#����iLL�CްF�T�p==�C���a��,�������ߘF�	Q��i[�I%��u�U��A������ǒ�Υ�U�7̙^�����E0/�VV'|D�#�i-�V��]Y9s��]��L�W̦���g�7��3�������Ԁ� �󎾾�9w��}����2�o�9:��b����{��4S�Q�@�wT&��#��ǂ�!!_�����-�Q�>��L���2�T�p��L�����8Uz��DZVP0#7������RBj\3-uE�h���T�L��er�j�����RW����/I��d4����!��B�
������Y�BX�޾��|�y�WoO�E��Rx(�R��h�����B��_!W�b���~�����4�O>�IK��T�5 F�����K���ZiY׸��_����{D[���b�-}�W�c�O0Q�z������b����o�{[��G��v��!�^[�Y���x���?��^%�ϋ$_��f|�������X��ݩ�0�������^a�q�ʹz�P���x
��Ά'��&��5!d�ywê��Y�(Rۜ����=B<�r��ӖlH��YXX��%�r����ÇA�"h�ֿ̝g^Y_EO��B%�R������U��a������a��|{�`G�>���f��؅h����ʑ(NGҍ��ؤ��!k��=�}�H>vp���s��?��[��m����Y���̼�>LS�¬j����0�XZ�'t�^�v{{S��^B�7����ٱ�߁=173���'��k���^�$��ҧ��0teaoo/:�U�)���]��r��B��:�5���d,�{q�"||���ՠ8�H<�y��� F���UU�r�d�-f�� 
��׶/��!T���(ZW"T��*~i�ͯk)\�ZHP(Oi��Ä�pqez��x_K)�Eu��<US h��뾎��u�O{��m�!���>[����`�N+b!W�1
Q9YI{~�--������z�>����`=�:F����B�KoHM}t�/|Urzzi2G���s�r�9>��х[�< 2�@�	�|�ʿU�\b\��m���0O���!�����F�[���x@����$$��7�4/���QVT�]_]�z����Ã�p��_m�<<&|]AQ11�@j���)>!��D}z����dZ�Ԍ�n�.��U��_�E+�����j�S{4i��8��)��r2=����sú�XY[;����:p����B�@٧ L��}�L͹�蕮#j���6R�����ꪃ��j~>��ڥ�z4U��x������M����b������d�i��l~mm-�6#>�B%i��X���"���X�˶�F�~������:7+��!����)K@Ӓ����zK���jkf@��L�%�,�h}j�2>�������7&�=���I������p���'Y��s���cW�^^��݊��!��?d!a���^g��(�6|����;,llΧO��wܑ��N�d���@����\�duP�C4��A���?;2`o���	$��"��ΥW���G"���U�.�������n��\�n�
j���l
T;|I.7'g�Vh�6�F)ݒ���G��-���d|K�	���H�L;�`�%,����4���n' ���.�2,+����+�]�z�탵��rK�9tpSr�kɽ�m�JKc{E�hD��
�S�r)mK��a���� 6�:�{�qC�_��������	'|�p��$�������@h���V�������$Tܯ���h��q�m�P���
PM.-/��<_�ҡ�p�߇_������io�K���o5�}~�������"�V���g�>2�2q���1�"�Z�>��==��b� ���5b
z|�5Pr��f�W�}'r
�oXͧ����=Dbp8<3�#�����t(Y��0c�.f���S��`(�Qӵ��	�9�e+x�3"S߃�a�pʺA{Lǽ�����,:*���V�iuH$�P��W��W���7�*��g�7R� 	6<=m��FQ�$���zT�~/��q�GV����'|�z��-i1{vA��E�+�>����_W/ƴ��'	r�-�rs��$8Ip�����.οv�y���h�:kiу����e���R��R Ӣ���ihi/���)�*��o}�Q����k��E�ԭ��A��3���=ob�aZ�����=
.8:�?h��ZWWKs��I���އj���D� ��G(������@*m�K����uҎ��Z�Q���R�x�j>k<�͂u�ȼv
o����̴�ZTY�}_�{�t�~�T�p�nt;,s�c��zn$�^Ť�+=���h��� ����Z٘�`���/������ef����H�{^;���d 0�:��avVg�)KGO�Q�ƌm;<�d��W���t-k��_=haM�(&��9ዸjڎQ�Ge�9_�6�RH�T��ҳkY��Wo�����ԷwZ&+��׈�"���!���r��� �� ���`�Q�'��2T�>�<��p���{�!���7 ig��S�=ޚ�f�k�>��[f---����@�B�^��f����H&�<%�ϪV�������K�#�|��:�-��3Kњ�/[�7��.���ML:���N+Mh��e�_��^�`U�Ҳ��" ����F��~����41�k�w�.��>�x$���9��P6@d@�|�=A�]�>�'k
�6�~2��/�<sJpt�#����Vt��B���:a��P,��t��+�K�*�8+;;�+�Cb���؊vw+7�p(���R��������@)���}�hԹ���̣�x)���N>���w��^v���o[[�t�<X5����0�$;p�ܯ�B�hl��X�ϣ)f��܃''�j�a�@BJz��A�&��؏v���߳ �S%�!�_����d�v}��T�'�~�nt�]Ntt�oޤ��v,z���La�=�Hh�xz�bGZČ/laPEK��B���#�!(X ���Dlrr���벲2Q��[�Cs��C?��,�O�1A�����>��o �ޮ?p|ޞP$v�'"W'�W�|�`����7	�VV�z�4�J�[��,�Qŷ��P2�r�@3P`/עS�w��~Nq1�֧ͩ��������R�T������}���̷�[ZVv�w���|�8��709�{qvL�#��]�I�!��0g��j���m����g=�����F���#��Ň�;9��Yε'�_�엃ֈ�?���*)��^�ň
;@3����YY�^R^hn��<ֆ��}��.e����폏w�}��zk����|ih��?���J�������`�� |r22Z�O�n;M�%���҉�cs�\��.ڂT?r��m}w4�� ��x�;^^���0��&NCS�� �Z7~;�e�dx��Iw��Qy���3	�˥tx|�:��.�R�����O�	���g�-<�\�'5�<��[�>z��
,��^s�o�3N_ ������}�t�!x�^z� �s�t�gCP0��Sl��A7�rπ]?�M�:nѡZ�F�u���)���"sDD��̶��u�K֟悆����A+����(�����ZF���odd9@ I�k��Ac�E�����[�Ym�\wC���7ǋZ�O��<�U��Խvt,��b�-ECCs0i^��N'Kv�VRRjs�8��\fOV .�p�Y�Ύ�:�~y��f���eff�י�0h��p���b�144������D��gq����m�hs*��g�qL ;U���pC�����2��P'=����^�0G�:����`f2�2	XB��d���f�Z�;��q[�n��S5?��͞6����E�ꑀ�������baK���[��_>0Cj�)���N�G�����]����rm�)3a���U�����0�:���ܚ�X ��M`b���|�f%�]��k�M�o��@P̷g��,cٗ$(��ttttd��I�Z +y�9P�
j��9l!�yyYXc�CR�Qư��dǑ=DX�g5�<OY�47�U6�=vq<ǚ��W6���需����u�E��?w��u<G"Օ��~����*�լ�䂿C1򤤤�B�v�s6�.�-�:ȼLJ��g�����s��K(��j�&�'��p���Kl�k$D���m�45�d�pexh���G���^�⠠߇���6'��8IIH������L{#��y% m��~���? �Ru����OZa��̶�' J��v�-�&w�(�o˭Ń�;����; a��v�ޜ(i��J�U�K��:�e ���:͞Y��r��7�s}�d`���H�+�j^i)G���]�,����^Nr�O�-Y@Hz��lq�r	����2!�`�o�� t|�m)�S�r$�!�((���o��֤���x����`3h��	����(������"��A+h�	����?5�������U�윜0CuPb��u �)��~�%��vxxz�#p�����T D��;�����M赭w�V���)Vg���椧��F)j���D�@<\�FK���g�HcY�|k*��_��0c���s.x�f��̄[�6�������љ 7 l��g) ��p�i��:V��żA��Ã��<FCT�nC��������k�@�Y!����j�T��uh@J�[*ٻNL�_�"?� �N{_`��:�f��1*Z�J�򞕮v{u -���ߕ'��1QiK��kL��o���׍'��[;��^�֓�������J��̜A��F���l� �U�XUVaU��)2?ʴ��@(	�$��H����7�t��>��[ �������f�I���5� �������Y���  ��'Ew�Lb4V'�7dkT�$�"��ډ<����A�LA_�Wg�S�tOFU���"�+���&E�6�31�SQ�2�"����h�������_������_����V����|�A+�i�<�Xf9ť��b�ϩ��%X3c���0^�/�]�FzW�^����E�վw�ǉt��U1��6�c�'o���R�������ק������#��r詯�;]ϛ,��#dր&�*Jf����x+n���"���wR)Ҩ,��� ����2���B�.@O��[򞧆�&Y�����L������h��� ��ʛVWO��ee*��[4��2�-��$�q��**Q �p�?����ܒ��c��mw��2��h�7~���6YfH9�_1ߜ,�_����W:�ui���}"�:5��O8�^�����J8!J����Z_[{
�(	��1쎎C܀�9U�ƽ魙����C9��u1B�Q�vwGܽ����G�|�_��:�'b���s���?��B:t�_m�`YrəЉHU��AV���D�����������I=d�.���9%%Ja���B��ۛr������
�J� ��o���H[[3Rx�&�(�ܼ<vx���N��auci눛��zfdbj�����'h��JCH��X�=�Pf����^�����U���w�򐄜k`�Z�d}ss	r�AiR��ɘ��A	���3g�H������jK��s��|TG\m���@��+��aB��al4��|v�ܣ����~��;W�-��#�8&��h�A��Oo����M�MD����)
���Y�r�0q�e�����\�М��1�h����@�B�¶���_O�k��K�jj�喼}P��C�
Y�ШH������NJc�W1\�����'�����;�D��ݽs'�^}}u��3��	9",_�f',��Ó-N�lH
`�����\��8�����+����G�$ ������E�	�2H��j���{����?K�67{&�����w�3ib&N'�dA(y?|��II���D�qo��<<��a_��o�+�:�- ��?���o��̨�k���&���Ǌ:d���wM����>��D[�O}ßw0��n՟��su���O���!�Y�@NG|'qC��k�B')P����
�İ�S�d���92---X~-$ �]q�(�Š�c�:���k$2��v�(E��M�$C-�15��}��_⃶����|z�6�T�vjQ��铴�NBg�D �������=���ľ�J�|�:&t��	߀��9��r*G�9�Z�v����Z���${���BShD���<�ł;���Ɉ�nmYAs��ݤ�0���E����቉��WnHI���śvש2�ȅ��;-�Bv� ��|�"ũ�/'�)�ݛ�AL�7"e�q7?<+ЪR$��Je�yZ�}�����P�ʩr��[8M�8�,"�>9/���G�v�jpppWggܡ��d�P5f���g0z��_\A}�B
Η������~%9�WI�Zc�xG�������]x3C�֘��{4��b,�"�-�kz��Vu�-�);I��o\�t�m���|b���3���]����u����:O���Diii��f�&��S ���F�S���$�/$(hu��S7��~uJ�B��|���ũpͬ�T���C\��K����3_��B�0-��i�~Ǭ��	��Oiz�>���d�w;��P��S`�������LPZ�l�G����<�� �λ�#��D��dl�'m�'PD����bfD!	�&&�Г#��мdu�b��Z�� ���q9���c�b!�Б9��h��ƟzB�S	�����i咆;#h�ʡ���O;I�չ@���@��4Y�^�F���1յ�~��}V�/���}�S�--�1�c-��&0� ӣ�;�9hN�6)�]�mA�va*��G��DL�8�1�}��ނ��ڦ��A�m�s�H�����qu^ ε{�hr�?�����t���݇��N�F�^���}�)�ݼ�6t�߾B�nK�Η{��v�!��v�82���7�{d
�q���p�&���b}�#"���.���xc͗��)���|BDOG���s��=���>����_~m������Bq�ZZ�P��6`gg���2xw�F�0d
�h \G1��SXB{)����iC	}Q���T���֛������YX��h���^��?����z�x%<�>C�@�'x����BaՓ�پ�~oKp��Mg������Ɵ�@���~\f�m�kd׺������`��?�<��{��j��~� ��W��_�y�����o�����v'��U���3�1ߙc�1�{�V�П�I����!�s���ٕ>~lVU��9�+pd��ln�8kY��l��K陂� ~p����D��E��pݾ=1�:�|����fӫ�����y�,�I�lb��B&�5��N�b���x��0X�O,��[�(ɵ;&�\I?�vE���k&]!���G��;m�>�߳q�}�wg�#�x��O�ʫ{0XO��]߭��l�C64�	�GGG����U4Xʄk���������v��҃iSKK˭���	G/��砷���4�a�K� 	��%m-��8�o,��;�����(��EKP�u��hҳ��n�2M���6�	|�k��=./���i�:�ʺuFp�2��(eA�H	�2@#*R��PCsPGAMJ(jD��^�c ��%H	�k�0���O������ګ<�y�9qR���3�4e������In�[������t��3��,�r���[ܡ�����X-Ou��*RAdo^O̐��|�g�i�[]�F�M��e91�/�&ۨ_�e��i�b��ҞlhH&�����Fnb���,v��rOT����x@k�c'N�xf�`��1m>n�5ǩ+C�h�H2	r�_6�+�����{���S�377�o�9�z���e ��J�5��omG���g���>9LZ��G� "���h�Kz��g���C����Ӄ�]�������l4Q5����prɧS���{�w��F��|I���p��`[{�ڧ��w�� @g��=�3t����A#�W}b��������a�(B೮������\��a���R����L�A�	5�:�0�H܌ HV�4het����o�?	�Z�Cf��T�<{ �ī����.�S�kq���:��L�n"�g�_�ڊ����2�ƙC��>���Vo\y��C�/�f~���
�<�����%��@��IQڠf�`�����6���U��<
��_]��������4嘿��m��UN��3 6=��E�@�M���o��\Y��/�"�%QL-�=���w�����]���_Ƌ��x���X,�k�~_ۿح*���-���=���T���Ǝ���o�����\>��2~�h���<yʞ��{��$�^G�~�ZF�Q!9���n��rT�*dj�)*���8�8�|J��nUz����_������E^sK�
�%��J��2�-q�x囩ja� t��턽�6?���O{��?g<�FИȅd����X�C����S�x�G��(��J���S��8)�/.�����{b��������⸙a���U�]�
S<ت`~�����7$H����_L]m��"?��O�D�6�������P�%r���0~p3p�@�����
�yG�֧���y�5�b���Y���Fh��7��O�!��UV���%��v�� N�=�:ז�?�%<~��P�O�(���0Rt��? 6$S=b�'p��`d�1�%�"8�U;�	>t�p�w�y�i<�h?�Z�yhs�=�q�`��0��J;���G�J:=����.j�)aT�0+
�~�]Ay��#���ڡ��	��o�q���U}�E��P_��e�0�{�}�S�E0$ݭE]n�)[W��?͌��V�IZ�Mt�v���S̛����q~s�ů�١���z��ez!�J�@a;`��J.����a���F�Y�E0,r$����Dz/�"ܨ��	�����2���ؤq�#m��Y8��f�x�+��rC�9�s���v����]��:6�����l;]&�&���x��f���B��?��m��O��gb�Ѐ�*o�!죮{]6�5y���H[��}�*����z4�[�VW��u8��܂��ҙ���f�k�:�<��N(�蔦z�{sa��>���9�Ͳ�U�
�_�7����et��<���YE���_rv!�C꒞���bJ��E�gV�CL��}r"�%��|�g��ϵ!{�o)ܒh4+��f���k �����#����u��ȶ�>�&���N������0�<l�'-l�z���G/�2� ��iX-�
 <Ԩ��2QD��K���;�W̹Ek�dZ��~$��_����n�4��8� ���Z��v���O���A(;)>��]y=��@�Н��(bP��޷���L��!�R�q}��2m���%�,n*���<�����B��=_2����#��fe��k�M�xv#V��G!�߼��0G^<�����X G�⒒�*!ETB�f�Y�U����9^Bs���\\���mB�9��]������U���@i��®MA�H���t?'�lv��F�S%YX cO�F�����h��	r�U�FZ�E�܆���	�ҁ)H.T�)�7=��WD���<x����y�Mbܵ�L~��\K�S�\gҢ���^���(���l��z�K ��{�
i6װ�O��]���ү�Y_7��
X�!lhwm9���>��,��Y�C5X�b���KP����2����$�E���2v��r���[��3��n�� Z�Y�h�����^�/�f
�p�1l�EY�Zj���0͹^�^�Kā�#(��V���e�-<z.E���[,oU�4��x!e�s��{�"������ٍ��k�d��Jq�Q���]?�r���S#*��b��}��~9��X��J<cA�S5��v�4C���C�t4���D��R������ʏAd���Ij���Yև�g��E�R���ߊ��ǣ� �)�>�� �~=e|ۇV��b���h��~�U�����G��wU�<�S������H-�Յ:h�o�s��������po����«��/r#2�蚩_~p���dj�L�F���?�@��kl���p��T!�|����a��m����fx^��H�U<eee\K�?Z�~�i����ӆ���f0��{ZŤ�8�b��P�贌↠3�$��ꫜ��=��!�ޱ��,A�'�:1�S�����+wq���]������Ėf�N7 Az7<�􏲸~G���p��Pq=����ք!��AX	�U�F�2u�|H��}���{(�X[b,LLL�KƳża[��:��\�\��VJ<Rs�Ԟ�cXh�έ�Z���|��ß(�'��ʴ���MU6`!8�4�H�����x�?�=�4�d�юԢ��4eď��<�ܥ�G�U��R�://o�Bc	x�u���a2#�i�-7�$��o�����3������ۢ��i�G1��Z�	_����7�z=E�w���G6?���-؍w����"��P��'���tTMN��a����ŏ�|����x�Gss0^^�����`5.��O�
#��d =-�b�:�}^�z-����Cڨ���)K>#�XؕT^^�ȼ�4�{����3J��Sq�W,�V�wu����^�Z�7�Dr�D�yTM)��w�;!駲]��>�Q�alΎ�xd�IFS���� 2���@�,�g��)5�����.�����&�g���>Y�N��0G<����1��6T���E��kx8p�sf�}n��
�Ё�����>�U#ظ0�Y��u%��M[�2	M
�F�zG*J%X�v�@�{��4Ӳ����G���3;� ���rQ���ӳ���2f����H��R��6�,M&�'˺~U.}���P��=ҝ�8\ ��i��W��3J� ��W:C���շ�]WWz��T����w�N��M�ht�k�'�#�%��,��b� �D�qQ�����}���Oyzz�J&˿��Gg1ۓGl%��j�g���g�lW��Y8��1r<���a*Q�ť��� ��Tۻ([2
?���F�����4$$Be�w/�#���d�<ҳ�]�p�&���٩7��A��c��X:M*�����#�P�Z�s ˡL?S+�s_{��K���a%�7�<�_.�F���ǟ�g �$�7zg+���M����졨ȁ�������{�pq��/���j@?Y�
��Py---�!%}����`�fY��DYb>|g����[�޾}XP�<Q4��&�)��g�W��_��"_��|�Y�ˮ/�z��=32����M��v�׷h/����EU�`)��x��
dz���{(�H����j,4��A亹_�[<U�}�I�5��7���~���@�ҔE~D�C��I��������M[��	�����ڸI�I���V���A�K�N?�&< 
m��b�S�� �/b�Y�����h�{�Ź��U�Ta-o(i*��(X��I�_h��f�S ��@a�ǈ���r��9�&��W��$�R������#in�ǁнiV�� ��t̋9vwkD����K��D�Y����i���?���.��8�a
D��9�)2`�l@2���z�F��? �dl�|�,1*j#�3[ف�;�)/���gR�1�(��dj���HBR" $^��d��퉤��e2t�(����=�5�zjRϥ��n5j�Qk��(ٝDp��<F��Rٜ��E4o��k�Je�E�h�TY��]���G_��"jW-��؆�׶	�)]YY�0dt��*��W�禒{�E�>V�R�|O9@DKa������<T��~�|3�U�ht���p���i��7�������#�տ=!��fK!Ϭ��g_z��Q$�iFF� ޒ�]�@X�G�r[e1����?�67�!���|�\7�k.����,!���Vh)��������;�?dQƙ�]Oo ��g
J��H�\�Et���!ݮ���[�z��e��7��>�rM!ͯ�T�����ݭr��l�GKmy	��)轮����(Q:��4U'� �;�Z��oV�O��x�(gk���3�HM�Tp�;kGA��ӹ�?v,i�����o{|���#�O�<yB�r�����gӲ}��/,��'e���X�N2�����>��L�9��N"�+������a 9�a��Xc�� 5b����Ϊ��x���������l�M�N2mkn�]�t�byNs��f�۶궤�n��+v��g��_/% r}G�d�U�"��+���);Acj*���`��Yf�L*(_�-D�8F@!wh��E ��!��gin�z�v@-Rw��T:!v���b=��R苋�1�U ������0W����S�W�#9>����7h��瑄m$t|�0�Ll�CG�e�=�|�pŤ��>�����m!�:+�'5��?���Y�\�:�h齪�è� ���a���V���L2[��9� ��v�{���Y��lrHE/���%V�zO
���F&b�gݐ�΋�
4�:�8as��_sb��v�.?��oJX�I�hI�s6�S��3-�p~��4,ϩ��#0/�԰��܆�����N�֣�a&>�])�O���o�47A˙;�=EG�Qv��f���##�ݭ3}��j�m}�퍪��)��k�T3|��lۺ�V�c��?�׉�|���l�i�6��Ar����K�Q�<�:EX��I�a��T�$���\Y��Sx����1勯��̆_�	�ݰ]E��O+�,4�kN���8�����,��  p����gNv��	ĩ�ъ��>�ғ=$0�[�v_�H;��*\	��۷ov mE5<� ,����d4:��D�8�Z�P��1Xr�S�	X�_ʖ��>w�y���w��V��eo{z؟�
Uǎ�ߏ���G�jE �%�fV�4ϋ�q�8a1����S����5�^�w:...ZN���q�v�W�>��~�+݊�@����}��'���l`e5p����-I��:����h�{��7f>� ��k�2�x��ӓ{�1)��4��--��g%%%H�RN�.ćE�N?7��y
�&��pd{��m3z��ùLK����-��P�M���Ů
yt`�Q�f/q�����g�U��x���fy�aʚ���H�xh�(�o�//�֗�p�O�P-u�Β)����g��ñ.@��*��L��h�sصQ���r� ,8��Fh8�1�У'�&�����n�A@��x�Z��r Q�I�%������%j��(f^�ɑY{����m��إOĆ�Xw>?��%)>?K�*�/�KܟURgB\|��x�o�D���sh�|���&�)C��=�*�	`��涎C���R%�b�t[�)��"r��6��w~�˫}�/ο|�N8p�,!h#�$2�r���L�	��bw�5�)\X�=P�k���;��fԤ�ny,��|��j���m^���ڬ|���y2�6f����Xq���K��*a�pl d��A~ CGP��W�.��p����-�bex�]��_+d��S��V�f�� l��GZ�lzTy�cv���y��5�t����m��^.MV� ������K&�tT�m�7Eۯ���f��{ �y"�'�ٜ���� �O�u�#�3��<P,�muܝX�ϒ��d7���Fg@�$�/t-�ba�߿�=g���_�Y�H���'�Ģ\�Ï"ob�_]��	lr����١���+�(���j�w:+�u�{�	rT�D'7�>�"���*{��wD{Dn/�M��EC����e&?���=�c�s\3ͪcT�Ư�]<Iё��h_������a��}�?�Q�����M򦒕�1���H,���B{��,S����6��KcC�|�'ᕈ�N%b$!@;��D̶��;�=�|�{DԞ��6��5q�لf�t�Q�����z`cnͪ]v}��kw%!	��)�z����YR��#�2�vA�P�zF �,}x&a��u(}ϖ��#�Z���do��C�����l�����f���$e3�4��a�B��Y{ƛ�H���,��&��#�@�	I/b�������R�Xg$����
-�1�2��� ��胐�2sKâ.E��T���������=I��D3��7@bA�g�G2�t��j֤O��W��W-�6HA��
��ZƛbL����/m���"�:��"v�͎[N�~J��	+�x�Ow�{�ݭ(Һ�>�o�����y��'����4"�h$AFGA�q&V����0,oW}���9�r_W�{���W<���+���-	����׽ӭ��{���#|T�?I�Y�Y^��I�U���&B�D���,�u}�;�Q"�e��\�蝭.Ao�m�r�����O42/�jE��S�b)Y ���<���5XX��D��be���m؀Ǚ�
h)�i���NN{�?b`���=�`��5}���:1_���}_�����#}�� ���ߩG�I�$���oQ���(x���)�ڵR�Q(s���(:�����gYZ�6*�-�<���@�ik�1:�
&Z\�ê������������Cgшmz�n�p>�ΦY5�S�#�|io'���"+9�|�4�Na_䴠G�\�{�}Mviv��f�"�*m��#O+L4Ƌ��@66#��Ҷ.�[�ob]����e������F,yQ�5����4��)�Y'�!R��2.Ģ�%�ooO�'Yy�R�)ɟ��W@�Հk�����_��xq��,DP���̮�;��wD�KM�O�-���s��Q��׮��O\4p�Pq�|��w�À��S��Iv���<krbz��(R��y$г,�� �^j�`ת�?DL�%I�l�E$#an���e�x���R?��r�)>�t���r(�,�O�d�e��~8��R�U2%۝��}h���V������V����GHS�|�� 6X��Pp��r�¶w��M�x$:K���GE0}����	Pnc���zm���a8���]�ңQ�
i���{]D�[�yy������h�����q�=.H�E�;R�D�*��S|�RЙ�i��YD�:�L���#	�_Z�1��L�໎��8inn�NQ���e��nzg�Y�O�B�@|h�K�sA_$1�/�����"��rrUr-^�t��L$�+�JN�D g�E�:)f�?��]���Xj�g�'^[�>� �Mq��%��_N�=�o[�m�Z}"���>D"��~L��w����.���[��;�zF�}��ā�0�(��4ˠ**"4���"���1��z̍mF�f�1Ty���糲H��I���?L5N�����+��ecTּ@^H����,L29X�N�KM�UI��]�^
�fԣ�?�=��z��d�d�n�MMΆ�������$����)-���%+w����Ut��&��d���zOO4tfi]�����:-4Y4�h�B�@��u��b����y>hH3��Q ��������J#��؍Y��O#�`��8wU���ȷ�9J�Q�����a�>�EI|���ʐ���9#�(�;��&��%:�wt�M�[��b�y�ۥʹ��X��F����q�P�z��������SR2R�Y�7�������rjz�����&�K0����w8�Iq�2��c� ���~�k,y���^���?P��O�;𖕌����|�Y�v��޻�/�v�O;��}7+�u����S�F��Qw�N��<�U�j�r8�y���ƌ��*doR����cV�yi�=�A_��w�:x��Nw�w�����[�^<��~���O=.����bQZ#{��h�km��������.�����Z=5]�b������;�(�c̿���7���-hw��3wǍR��/ymW�kږ�(F\���~-ųkW��n�d�����F;�)�O+H'�Tg�{��4�iܫ��߫��(�{�����o�^�p��ݝ������(;S��(�齨���U����}(rp�,�]�0r�Z#E��~���\�T��,�A���M����VW�F�����FN�2�������I~wZ������w�;�Ez=��;�K89��1�"�b�g�O�a�+y�yy�������Y���ɳFH��տ����,�Ą�������	�(�T>B᪼�E��a���s¢�V���v:d�ԃ/F�T-w�ro��ʗ"J��1�غ8�mzuΗ�F�d�Nj)Vhs�Q	���?���*��Z��].5"S��T.�\���EJ�N��^p�F�R�ږӟ�0�tW�H'w*N��ݺ񹮼�t}GH�`�'�N�,�AY5�?~(�;�5��\@8# *�A�w�ϖ���]l+��m�H�¾�C���s �P������%�L�ެ��G���Ue�k�,>P/���v]���"��.�[��e���Z۪�MEe�B!1�F���R��*���*�����L����O��h�^�5�Sd��s�͵��ז�Z�@(��|`o�*��u�S�F��0�]�v�Oi�NQ�C{{WI_�֊}ȌZ��e��6w%~!)��E����A�е�'� ��N�)F]��x|�IYq�z�	ˈ@3��ڹ%��ܘ|�:;s�%]#.:x^��hiK^�;�h͝c�sX�E��!��9p��].���T]3���ޱ�\���s�LJ!Ҕ�$�.�*��i��i�<��������5��M��x �a��jq��2�5#Mf��W&�;8jAd?e�����������fwM�� �2l=���QUe���Hi�p�̟-!�׸�݁��3rhG��y�k�u��[��j2�����~/n ��Vv�[E�Ί�n�bV� ��[+��n<�%5p2���K�����q� �g���f�KR�{ī����qݠr�)̂��S���E��F_�S�m(+���Ad7n���J)��ua�<ZU�^3�"�qA�#R�fR�7vͮmu�ⲟ�6,�����>b0�m�2m�B�W��\�PM�kFG�j,��p�����VnfG�I%K�ؐ�	p�K�L�c߭�?�,�k�]����x*e��e��5_|��oж�E	�X���܋�;{T�uN�oހI���h�eC���6𤥓pǮ�C�DbQ�5oGi�x��'Ba�.�YjF\:Y������w�O�m��k�%�YF�]s��2�$�aQiCP� a-�f=1�"hGE|Y�#�R�X)[�`ϓөg��c=	LAK��Ɔ˜)���Le4 �9���-Sp�< `uƳϽK��X<-�#+~X��3p�tD��7�'$'�����>�4��p�WȂ�+i�igdM"X���+5i���?.~���p)낸��#�
�αr�N��+��m��X��Ű�a���z��4�?���4+5�\��:)g��c�?2�X��?PK   ���X�ة� � /   images/4cb229e9-cddc-4c52-860a-b86ee61c7037.png4Zct]]�Mnl'76۶��F�ƶm�qc�qc�N�_�o���>?�^{,̵�<gG*+J!������!�H��~�a``���_OF �̯�EUJ�f���LF\D����/�������zje ��} �,"
^K�v6:
6�q3:* �6�@|P��FED8a�K�AM鵷y
6�9�k�q˓��s4.�����{b�7�sR�������r�xm����	5���x=�$	VI��\Ҳ��L��6E����ZܘTIy�c��4n����bO�������'z�<�Q�w�ڹ�[�@��p���UܧJd��ʑ�T&���Ϝ�F�\�|��Q�Ώ�o��������M���NIg~�5-K�??�-����;��C�Y ʥ�W�8����xڋ��G�K)��Sq�U:	RBt�O���eP.��rΧ��3��nN�~�]�%���L����9g9~�@�a��z�Z,�'���[��"@�aW(5!��X���d����z�-3�c6�,��T������P+�);�0Bg��|a1�_`�@~���b����'�D<M��V 9����-��\��:�	Јh
Y�P�}��d��ƭ�;n�+[�Y�{��9�y8���Z�������^��lG�k�I���o�]W[N!p�]/�Ur>���I���,	� ��9v��/�^;)F� 1���u3�UT�_���#����������ڟ\��ܫ�8����͑�v�����{Mw�	�ם�㳹�qu�c�)`e��/6:Q���/zɮ���� L�p�<���,ב��v���G���ڹ!��G�'q����Z%Y��1�]��ޕ�r?�)��t-&��]�5���� r@��h�y)v�;�?r`�D46��U?�F��?"��hʧɲ�gl����bŲ������O� _� �ƣ�n�1�5��T�<���u����d�Bm��JGq5tj��Xl>�}3s ���ےB��<5O�e���HS�y?�>�-nw�n�2�S��~R�q���k��k�$	UT���n|�{;��5;�y��Ñg�
����,r�vc�ߠ�Cvχ��1�����ٸ=@Iĝ��Pb�.&a	ݫ�&���|��|�����6���P ��i����u04R��pM;��.*d"�T���b[�4Be�\`�G>���z��̓�����y~�:�h�Ϋ̅*�-��􄒈�S�u�Ɛ Ih[T�U%�w�+�'{~5p�?|��wv��Y��*�y�8���5�p�j�k��&x�i1�I'!"�C#��Q+M}�/�
Լ��js����a#3�]�+*i�4c%���
dLɱ�ط���[��Ϲ�QQ�z	��+w?�w�xyt-�if��ǆ�	�&CM2�Y�D�Z@�:�k+Z�F`�=�Y��Ώ��]�,�ޘj:,T.DVy���7���!AE=��u�D�&;���A������c����H�6L�T����f������}&�5:|��5��FF.����7z"c#�Q�vvfQ�}����W�g�"��q+�ϲ���[c������$.#��x��ސ���S6�jA�Qx	�@�rG"��R��{���S�U���x`���x���[�R��N�Qw�\�5Z�L�h>4
���/�%�x�7V�u� �,˝SFe���Å��� ���v���!|�-.�oE���?9]Պse� �\��찾�db�`̢|�M�A$�s�?O�	�gw���%�y��u�ʵ�s�ړ�1G/�f��?�q߮�#�OР����2�حg3V�!��`ȳ����tr*I+Hǰ��s�M��̮K�;8;f��:��u?��j^�q�F���'N-".���Z�o�`]|���s�Ƀ�F҄a�I�67��6d*�0
���r���5zT1�c&��~�B!O����L�`9h�SV�9'�T�<~��R��TEEERο)%ï�,
�������j�����j6���z�-lgK"�ڢ�"��n0��MV*�e�~/��yX\&����[���f��fQLLLL�Mr� mM� M��U�|����#O��8���~�E���{,ZbF�v���J�a��h9��6� )���v�X�b��w�!L�u?���Jn>]"��;���2���b�N�"����\#��w�:�M��?S��?�ɿl5��|�����.����cL��?b���D�E������E<�:��r{���,��H���50��^�XMC�����d�	�_#�����A���6a8r�Q��o�;ڒ�������l�ۆZ֖:p5^ȯ�\����Q8�az�0�+�c{m4��[æg�|W��JYx�M_�.�j����s .�h5XK{��&��!�A��l�{P�Q�'@D���ڟ�y��ّ��|������q��n�d���c���#����i��0�9ԅM��n�-NI:�d$I���ta��̽���$6�<F����@Ny&�=�D���f�������z\��'@�&�Bl�c�RC)�h�����;t4T��]�1 ��6�4 
���P%&5:�L�%x�٩}�UUltD�+]�&�9�7��	I��e���*g��kb�4�'�=N-_1�/�Iqt���)��B�7/[�T�/���N�����ҭ����or�u;�Hs��p1	���&��t[k���F���G?�K���Mi;u(2[<�zg�T+c���*�4�z���J���*TԶ_��Y���^��=��D��1@����NMK
V���]S���,u&��qÅ�^�4��m?M�5�չ����&�|��O�>@�r�����72��]k��y�#�����+�W���&.�O�����,C�8o�D��Y*A�ê>t�Y8G��^�B���N�Iؿ+pq*���Dw���2��aH�hhp��9�ξQE�����>�|B��>����>���[�ya�����;84�lM����$����J%}��$-
+Ga!_��@wI^��IVlF�$"W8�Q$�I�}��pJw�M!��?�YU]a�/������W_8��苙���ҰP�N�6/z�he�������(�*�%�"Nv��R�����@�&��݄��Q�Y}��.ܗIʌ0��}�����W�x����#o���X0-�>����F�~��;�8"P<KV�)�"I4E7	�
��+4�r �M���TBr5�g͎���U����Q�Y&�g�-�:�3�9���K�^�4,p"��*6�J2[�0��e""-�!&^�\��6�� �eb��r�Y@�\��l��C���}a5"�Z�ʎaE@�KL��M �������F�t2�:�pA{����pRI0�$�h$�Y �Kd�K쥮�������DI��AQN�T�v���ɜ�R��׀H�M��/�PW�זv��D�]�Ѱ��,�+���I��T��u�):��de=�h�H��}�(���qK�h�!���w)��Io�C����s#���q+l���$	�~@�0�r�nt��{O��6�S�L�^���"��<�Vj�����F���<|�^ry��p����|��P�0;�1��*6�]��Nl`���Ѐ2ҝ���L��'.��B���oo0�dk��l���+p��m��d|	�ߢ���n��-/����=����?���W�����O���!cn��1��~�nڰ[M�@ 6�<\l��U�~�ol�D-��cZ-?e(ANaŒ8G���w^nmK,?֨����z^/��V����.`���VZmǦ�Ă�k-�d��g"�uڄ�������jLH���� �<�|^W�~R���V|�H��+��)�8,L߫v����t�*�o90h���M�G�/nޣX�7�;'��n�{D�n���F����9�A���ōy�n剌������o��]���3�O]+S׺�U5����}��G���2·�n�н6�`F�o��4m6K�l�
U��	��!~����%C��L�@I0��ﴸ@�-4���l�WO�b�����>#�p1	l�7�T�aH߆Au��}0�	W�-���N��%SB]l��6].g�}o��j�+���5-�s���^,��,�"K��{ c,�Nb��[�y���+4��~���h��Ԋv���#[��D����21$�n����8c�5�Q�ѥ������Ui�U��]�����g��3�` ��bEt�u��I����鶱����j��r�뽲��l�]|ɸ�8��4&]�s��:����_���/�yT�;��x9��!�0ZK��b���/�'�pEma�܁�E���y��Q���4)�����'��`�S<!_K�r�iz��G#��d�j[�������XG�p��l��e��|-�.�a�>��4�Ð�vޝ��_�o�������f�z۲�	��@���J��Zˏ�ƛ-�S}����\O�)�^��ndM�&��&믺��� ���.`�nz2t=�+�E��e��n��[{=.���5�wd�3�K�������»�4H�ۮ�X���1�:5t. �Ǡ�ş�m5Lgԟ1��`Iк�����p>���x� ����G�����^���d3��zI� �)���x��*g(Ģ�� ��"��&k������􆾶2u;et_r���8�D{7Ϸtl|(6���0CU��$�X��qfj��B,Ds���{<�I|a���\(&���4�=�j&�֗^6b����v3��u=�o���#���]d�1�������e8�Fa _���/I�wO��8�S�ߺ��?�_�Ϫ�l��Y�à@�_�m�K?�y8��yd�}��`ID���*�ϗg����n���B�jΙ�bD�����Z��R���)�k�*4 ʹ�>Ë� �$�S�4���tCL�5���y�S���ƺʌ/ �db���j��u[:�#��{���������s�q�[��b����R�3���܍����" �	��{)8�bp����
nr���������l*�*�h��`�;~�nX��o�f*�����AI��Q����.�i9?���oK��7�O
�Lh$���/;��q������:���>����zpF8��=�xC��{���uu0p6�|JIIa]�S��9S��X����r����,�H�Eҭ��0���Y�=� ���`���B��82�����7��	�|n���{kT<�N��3��l�PŻc��'��p�Dd�7%P�,G��~o�/����7�t��C$��:i�K�;<��
s����cw��26�h�ӵ�ï^e�l�Q��)����xG%����^
׫+9��A����8X>РA��7��R��8�������1��䴖���B�7k�]�Ͷ�-Xc��V�`W����/\r���z.{�_jGC|1^0��y�����9�eD��${!�Kat?���׹PB��0Vz�����t3���LB�s6R����;���o�?$��[��T�h�������E�ea���L�����p�\*.ǉ#�a��VM*�34@d���
GE3�H�&�mk�G�sL1�M}���8��"��G@0������C�Rʋ�n�_轤���~x�s�a1^gꭾ�^9���f�U̅���K���D�L�ewI9�k�;�e.�~���9^��#t�]��0ŷ^�
��������K�/L�455m��K���2��ٽ�����>�"i�<��nd�A�r�p���YXƕ��z�N���:���TR������V�o�H��|����D!<��Т �p�}�	����M�4�^����V�>�ߟnl�����w���+��5	�FD<֫���ȗZ�˵2�/������7�,ty����������� �ǐ4�d������Xu��ٖcBFΦ4�p��W�d=�+��={�����R_a���[g,���L��Mжo��(�6&�#JƼ]����i���b���_��-������@a�"��r$՛�Q}Ѱ������V��/>"dڶ6V����f��d��`csZY�ŶrA��5����yt����&�!��c�N|*�)#E�~6Q-�2DI���ݛ��j5b܂��H�.��q�1gLR���0�;/���ɀL���"�?,c�W�|� j��b�%o���W<��?�:.q��=n�~�� c*�r�D�q,�_�u�V8UֿX!*�؄;�7������U!��l:r[`�V�C�l�o�)\�K)��0�v�wi�y��	�Yv�]�}y���i@��d*:�ʐI͕.sb�#�h���%X�B՘�O�Ӝ��:�����G�)�|1,'�U�8�����N��:Z�$�����*N�A�i�C���*�gZb���C���@4���

�}f"��<��]��{���ֵF_AC=�H��ߚ�*z��(���[m�m�C���������9��d|��}��v��`bη]�L8j�s?��uy������ר��Ld�3�X���|N}���ÝLw�������p��siA@4��{�g�H��M׵�,l.�N��Ơ��[�7]��=)Sʯ��D�]�J5z=#E���b9��r����<%fZ)dF`��d�Z�C{��{�m/�p7�H)y��N �uW:��1֞@)�٥��z�"�����7��\�_�3l��w��"t��dG��ZK|(R�N��%%!9r%PA����-��������6�к��h���E����]UV�o>2Af,��p���."#`h����l���"�y��@S��*j��<��e�)�8��&Ȕ/R�{���jCmOG����?
�II{_ܜk&(�k*������`jh�iXG���l,��M�w�$�O���o��ttx��u>'8�M�����~�/��[y�6��v�E���&��t�f�����9F/����Z��{kD�~�f�JJ%��!��f	��=U���q����Xr@=���+�9��\�U�Lq�٨/h�+�G�~S��%��$�����.~U���X��,�)Q��$��UV��5��[f���쮐�-Z)�d�I���P��M���r;s���lv:��F��9,V�j�ֻ��]�������{Nl�D7e��{=_�F�y�3Z��޺�2Ԯ��X�9%�xT�մ9��tj��vE�$��~�wBq�\,6�5x�a8+bw��y�*�_��<M�� �X,'s$���;N=$�A`�W!鯁md� W}k!�g���ʑ�U�
�eC5+.R�8����T�'��ð��5��}h~V[x&`�:�i��>��e	x?���~챹��3r�O�"i2���`d'ʈ�^^��������a�1���f�[������n�OV�lۇ�0$|�p���T��/<'͑�2�w���Onfi���[w�سJZcG^
�#��>^B��z��'^K5����לG�RB���;#��21���/I���j��F
�y��|_�������s'�k�{�6 �Q��Y(�H(`����,LZ��4��J�1��?����s�^Y�+=��G���D��m�у�Q�Z`N:�R�5[��	zaT��+T�2G�S�� X�E�#�8���Y*�J�ac�
����8���G�a|����y~��K���T%h�#Ho{�ER�|�w��bL/��������9��h�(f��%� ��	��9Ŗ?�������6�?��-s�L2�E��f�	>�r��1�p��A�� ���	�j��ʼ�Ȼd��p�>��\��ǈ^�\}e�A���g/��/��~~���f���]a�=�-���	�1�87�x��p�a�E��~F4q� ����+C��_���#/�3qD�ԁH^��L�C��s��>���.{O�}�[9mJ�/��f�z'��떬�.aR�eh�AOD��by��αyp��(��
�S���u����_���'�2]\����l�*�>o���{�B&�z�b�ΜeBn�{�l�o����+���#~N�р�9�7�Oq��#�cLK��`Ez�U
H���'�"y�JcddtT��{�4t����0���Ip�"��O�_�'S)Z	�=uf1D��.�+���)�r����
	w�G*����*g�T�tw��x\T�rG	�Q(6�$�m�
�|zeT�����C!����`_�0��pN$��"�@>O�>��T��屼���T̘e�~���&����袂횰�Swn� �����K{y�n�%tlK�U��n8�����u�^�<>�-0{�!�!Nn��+�{m�g�S&U���k'|�����m�!��\1:g�LC�I�����5��
O�X�w4�F7�Z�]�C�|�[�� >jp	��,�Ң��Dh>ѿy|�@�k_:�F�Oy/�^?����8]��><C�oA=?nQ�����}	j"4������z��>7�
�ys�Q�+�I{w�������n~��z�3�}�L���M!t��h.1�?��������ƿ�n�������]�p��X���W�H=����u��2U��<��u�3L��ks4V0���+���Ԛ�'��f����۴T���h<��[e�}�������p����Ȥ��6>W��C^��ԑ�^�`�p�Ç��c�,"�U����ް�С}�XчըT��B�s�;`������=�c��ӧ��zi'�0"h9f�;��{�L�6]�U�����}Œ����?������F�<���Q(�F_ߎ �
�o(�<��-�>[aXV=�34�p���BFͣ!��Rs�\o����Z��z��zR�q3�}˿[;�[��)�����k0�M�l҇A�����{����t�o��g�jH�����N�m�[xN\��f�-�_�w�]��A�WN*u���L�e��Ó�r"O�9�[K��y?�k�FjK!�g�ѿ}��-5Ԧ�_�p@�����ݭ�t}���!3�ϼvk��B�8��F������Gb����U�a���w�����رR��},��'8�{��P5#�ft���5�:9¾��x� ��x��P�\q�����"Z6��F�;�R��n���{0�57�$�Ӟr�+��4Ň�y��`�d4��� �D�4�L"jz�H\dus�߼�P�<
�c����D�6�=����<t�D�a��L*���x�2W_����J}u�Ο	kab����4b�R�{�����z�!���`�}�K���ߜ+�3qR��UmE����H�EZ@OӞOe󀽚�R�e{�0"2�ze��*�K"4�j��x��|����,��5x�8C��"�����Qnu�]���h&6�U��m�
<^�vn�U��6�Q5��������	�f����	}al#��QM����f����M�)-�&j�B<�P�=�,���G;{#��:�HO�;��"ϯ�=���Ѡ:����Cϙ��ُFaI�)��t��Ym�qj~<���{�ӽ��y3���B�p�mk�G%z.5����!=$$,b�-d��e�����,�G�?=����I*�*`�*�*����J� mUs�.�@��x.���63;7$
z��*^�)��65��Nl:�j��a��m��rPJ;�svɆ@�9��U#�C��X���ڢ�m�������zG�+(���G� :4zM/Z�q[�i�W(ɡ"�ߙa�B����g6ח���C���H���b,��X���$�:��~�`���)[0���}�IA�H�{�d�27�VyybYp�°�_K#G��9	X�4�n�b��vgj=�EAMy#![�~�ZV��HJ%	H�"���.FMHv��;=e'Nő@o�x4�"JI��Y[E����Rp�z�E��(���J���]��H��T�l��NC�ҊZ�}��o�U��t�j`�k���s/��1Nd{O"��弧�J�y���޾�>*�W0�n��Y[re:8J�i���Kۻ1nI�׫�v�S]��uR��Іղ������[[/��OEU��ʰ[�FƧ"�D��P���*s�D[��B�l���}	g8��&E��� F߬�S���} �9�U¤F�����d��"D6:.���	0]�<|q�NZW�8�:���@�Ӑ �>kҶ�I�!s�o�8�^E�}��T��V��N>D����l��%�%��\�SP�(��y"P����u��d �g�+��o��(��|��A��WV�ڰ᷃�H�#1�q�$*/�"&��߾��d�>� ex�w�+jm�V������h�s���S��Cb��"��aA�v�,�ʒ�&�Q�f�K�Z���r���eW,{[,�&� �L��tkts���u2�H�l��'a^"���O�e$bh�y��z����#�r���%v�����J�sLFC� �+�|��98(?H���u�\B.�����N���+1I��_��&��A�6R�K�ʨ}`i����d���N�"D�uL�2��023�Z�a�h���=�B�iF��������� �fy����l>�ro7����h�:O��}{���>�q,v'��F�t��p�������,Y:�!c��Yga�tM�~6Y{ڌdF��j?�������z`֒�s�n`�5j.G�"�G���@>�Ó��KF:�J��u�f4���ϡ�F�>�]�v���Š�8�#� u���\��჉��q_r,bD&�v&7��.6�� B���.�e�N���g�'�<� �;O��%�qL��⟞t�-9��=�+X�n��pI�'��"1+�!��RS �oy�	�k�ޝ�ߝFs)�f
x;eo�QWw��Bq����C�!��^d|��b�*6�T���]◦T�KG�\`A�_�d[������,*�ތ)��-̒f��n�n��$�L#T�,�H{CK�O�- �P5�iE`�ᬾ
�TP��O�������n���G�(��
qIǱ��H�wC��_�;ϐE�4		�;[�9�˝'���+[��x����Xf�D���y�5�Tc�GrX��a�d�ϑ1>�z8����#�rH����М=|�̦ˇ_���� ��9Jħټ~?�Ġq��3D�-�өfbp�}�A���:P��i�=�v��\	~\�����p7���b$:��d�[箷 �%ʐ�ܮ��3]0�K����H�ĕ}{��Ps�P�Kn��2?df1�3����шT��
Z��w|3L!�X u�7���x��e�EN��T��9�Ŵ����AH:		�Ce�F{�������;�<�A��J�v�Y�\���n�|�+�׺�}	�.!�̇ëἳ��.E0��$A���'�_Pa�2ܭg��?>�
�й�i�ڻY�X�42��&}3�VDZ11�h

K,�8�CE������~5�`:n�o�$Cdj�-���3�	�!���Ա�/�C�z�z(`�d8��(Ig%���@jm�U�a<�;�0` 3�Ϡ5>QT˷n�a#h�S'� �Y�(�I���xKF�ЪX.u��*����̤@$��+(�K� ܵ�:��S�f0��!��t��p&�\���8���-��[hB�^�n���dC�(�\M3��l�FX�\3 ,5���*�2�;Nj,���p�ߑ���?��}�;�缀�f��,&�"��5 �M<l[�pΣ���Xب����E5����u��GΝ$YL��6��@���W�ʍ���s$5��NP�eޏ�ȅ��Q���Ytϟ �HN���o�>'��<�i:���d��?u4�`u���ko#) Ϝ��ʨw�n��´	��������#����CB�ӳ$BpH��uPW�0<h��t"��­�����,ǒ=��Q'�Ht��ۀ
J %,pY´t	����p�0#L��x��3�c��g\�|U�V�	lV��)�WD���L}<��0��#FƟj�R%�e&XmH%��U~�����s��kk�p7�ª�B���7䂄���A��T7;��HO �$K�<�*��d az�=d��چ;�E@�Re��܄�ǺbE�`%%�s�Cf�;�- d�
��a��<��G�3��;	B�4�-D���	��j�rE�V��wY�������ѯWZ ��6$`��h!�K���y�,�*�#�F�q�Cf}��4����b����V�E���x�X��nH,!�#�{u���{:�`���������4G�*���ī�w(��*��=�Я/� 2,�Q�͞<ee���}��sX�|��/S�3˵{�#{S����N=k������� "X��@���M��UNB�f���&��F8r�"�a���N�x�1P�aR�٬�qY:PX�X�(�]��vZ4%�Рz�����1��#�Ư-�C�]a���L�1xa�Q�W6`n"9	�� {�r�p�l$7����C�'�n0�TH��JG|�c2Oj���2š���FG_#�����\�K���^����|�҄�7@��}��=V�|>���fnm�2S� ]uY S���=�9E�+W��mr,��M��r_)^$V�
:�ˁZ���+Aݓ��G���w'l�5�N��NG�Q$���(N�[g��Nҍ�����+H�+լ���t�rzh�7�7]�+�Hٚp�p�*;��9�Ɖ������Y�qG}N��`�heq�������vŭH��@�(!�[���N��U����Tf~1n��#��
���v*�~���kb?�n�#aC�MPh�i��ō��k%o�Σ�/ꂄ�FW(C��@��}�I+C��~�#ubAn����}**!>T�[=I��r�+��EI1��i�c��C��5�"G����D0�`݀	�'NN�.Ͽ�FbOQ�8��$9qpb���:z^�	Y,1=TJ�s�o�����pb�� u��?�v�5�����ٞ�B�����$���X;A8�A#"|n�j/�ʯ�Q�+�u	��T��Z照E�(��^�\P\>j��F�%� �0Jى8[8���D�����m��Byh���,�4x��E������Vm��>�H�3&ռ_78\�
��]����� ��&N�i�ۖ"*��>D^a n[�<��4P����:g\�0l'��)��]�f�� �l�c7�&�X���<F�<>����DRʂ5���VhiՅ�CuZ�O:��~$&:)N�nr�:Wյ�j����M2/���'Q̙em�0O$�'z"Y !\��4 Ǭ��'\A��㑱-��`G5�RS�2����[��,׃�L�W���U*��ۓK2� �]�Y��f�Θ���u��@���kʱB��WE�&��p̐hn2!DW�K-�WZ�H�k�u ��f�����w��6��O57�F/�e��"R �+��΀�j�]�&n�H@ Thf6NP�O�X��w�w�sJ��KYe����T'�"zNA"�k,-�6v`eƉ�ȁI�pQYb@"$�Ql�<�������]XXǒ>�v�V�����	�=M��#:��j	�i��i/�r$��5��Z�{��'�к��.�u�, �����x�ca6!�0:b��Q�,�.9�Ƽ��*{��n�5r��CF4K+W!�e��:�(Vo~[���X��x�~X&�*� =�VI���p�����AQ!�uL~?Vy��ƞvX�<�no�¨D����w�ΗPN\�ه -��HE?H}�s@�]|�0���3�A��H	�qߛP���(3�qi	�b�M��M��>�;�I�:����R\*�]�����2��|��l�~e��-#֩��Tu4e���8�J�xN��mGִq1��|q@�V�>�_�-)��˞D��8���P��4��,T��Oy�i���B���N��B����/
M�z8+Hy���#я_�Δz�}m4�����F3�]�Ʋ��E�VQ8�άn�\s��s���JF{��芬529G�E�`?{�Sa��`F�D!�Ѫ�����/ i&�,�ZU�v�<��f����S=9e��K6���_���4���I���	D(�
�&�Cu�IP�X����E���OSz��@� �\�
��-�ʔ�9A8�guT�)R`�R:*�^b$7�%fD�άԼ�?�.�0�(C�hA�Ϳ`���4I����ZŨN#"Ii�e�S���\�hq���<��7K�0*��-W�|�؀�k�����j3rIڐj/cG:xO�,��`,O�\��6��YU#�¯'=x�u�G�����q(�jhSBI�hJ�2(�:�+�r�$�@���8y��r��c����^��!kR���J�	S,��d�m���]�X�mD�b���#JL<E�B2�6ȴ�+8���/�$�DMd�I�񒬼d8Dph i�~�:�1���	�H��{�Y7*V��uI?�"u�B"��4h{n�����"� ���M����Ȅ@Fki��,��L�\�N,.�2�R��K��u��S��:[i�O�a���h�x�qH�Y� k{"��C\��&�-�^؇<���_p2�-*z(�}��':aJk$Y�}ή�A9�/Ԋ=%� ��c{ W �IJ �I��-���x�8C	�h����b����0���)z!?3�LO�����Fç��ˉ$N_�M=%���TTCu�$��B8
g�N8IWi�p��X����jy�@V��'� �8�L�ʁ��Iq�i���%��q�"B�E�씹]�T#��זXf�<���;cq2�VRLp3U!�EYCj)�U���K���a�X��[�#�)�\��E3��I )8����{��^Pf�1c]=}�ݹ(8g$�U�=� �������{�̮�+<��6T9���;*wmf�����?"6,aa�dk~����e�&C
>�0��Z���o�M�y�%�H�d���V�0A-�̹#C5I8���? m���23w����[go�=u�pc���~N���y�C)���M�������6~@�&��*�_��Љ�����̿bn�hK�M   p�P��_1�s&�*tAK��;�%xJo\Ir�s��n}6<ҧ�j������H�ԲK�(��k�����R�
X*�!�^˭)��@���ɸV���A�<	Q��c��j�B��G�={4,3��<��o�TΒ���~]���ַ��������� �89^XG(���:vNbb!ºr��Z���Pn}����w��xUz	j`D�T� �XQ"��T:�Y}�_�=D���&��޻��񳼪r�4so����zweuY��'�b醙j,dn�b�l��F��|��zZ	ъ��X��94����ɘj&����C�elRZ��ct�b��}�G���[O,_�!���,����p8+�峱1F�PJ�fJ��1�������Oe ֞9�� �|`//�Ѵ�9�Z�ʶ�hGU>��m+l�h	^����9�,=�aU��3��)�6d'4{��`$�ݎ���8wX��;{o�Y^,�����?�R){�He���WB��) ˵B�{����~M�Djk����ԗ"g;jL�V�z�֑�i#���'�[������u� 0-Aɑ+Hb��� ����ѳD�WWߩ~�J��S��gNMʼ*�xh���V�$��eH�[�`����%_X<�Q���1��ǝ��e�S��
���� ã����)�)�f�/�ή<���J���UHz���LBj�$8����xT��v�өf�^W���4�%��G�f����T\�2Ѓ����۹��$�/`�w'YN1ezE��{��QJ{����𓛔��-2d��bG�!%��V��'��c���-R��.�IۧwC��J[���?�� K�8"���(�T<�}!�)ؓL�=�_������I/�� ����2pt����*1PJN	G���Z�q�ߩ�kv�m�o����v�J+5kj[�AQ*	�X�Ҁ1�b�?6E��L��)ƌ`6c��D)<@�+(F����^U����"�7mZ���M�� n=}I['�
�d���B�N��>1����z�%W˱������V��Mc}�����67r�D^j?>:����9@�v-��bf���mj��՛��g�k�����@�$���ڑ��h���^i���X�<�r*i�5��"��M�w���+���*+�Ý���)@ێ�?����ea$3]zC�}���h	������0������k��ջ��� �D}�@]
Ji�
�G�y�m��8VZZ�
v�",�r�"d�u�Bu3 ]N��B@���U��p��� s*����l�>��WQgU^}ĖB�:�v�)���.��yW0�n7�)��E�� � 5@ʿ��4v`�����2���Dp����� ��F�IƧPX[I�����x�dl�lA�,��U�(«i����A���̳,+5��9dW
�E�P�EP�U�WĈ;D)��l,��nS�EX}��aJ�ZJ��Tc�����\K`�3>HD�@��E����Ɂ�^)D����x!Zm���q�𞝈r8 �����B�nP�Z����,�I"��� I���U��<���N!KqB���SY�������� @��6<���E�� ��^�����VxM@�G�jq��9�āW}�{���,Yf�Vd{4X]ь;"
T�\�(*E���?-�@�s~�,V�����,9mGAn&��(�UEIY�����Y�vfԒ4
�|��oƅ����eIb8H��¢	�p�0����`�ZqKEoiƴ(#�[�P��ϗ��e��A���.� dʲz�����፞�3�%G����r�gǬ��bh�yt8�R���F�V<�
�@���En���Hĳ0�����Ywb�b��GMn5p�RC��dd4�Y��$B��rq.|n�K�/�2�
�� �8Y5��"�lV��d��{�s�B�0x>�� C�,a��K���1����
�����E��IEH_Nzg���.����b7�5f|�?m�^��n�d��b����W��q�v�(�Ω���1�V(�^;Y;bccQ%�@�u�fW�T;�v~O!��*^�lD1���!�TJ�~�� ��摗uN9 �+
^)�-��B8�S��T�0�����8��6SU�;y芟5!�a؝.x��@S�QV��L�-"
�

Ir	؜�,E�\N�șR�^r���Q,֤�JJ%,Ui`�8���
fX=�.� VMi�Ç���w�m1h�aܰ����1���84QB�Chz�c��Ŵ���K�GBl|~�%�� wUv��7�_v`���3U� �a@��E�
��,4���)UY��[�%������%���w۟�S�F4��d�1��w/~>�°&!ʯ�)�y/��T�W$��!�;��l�����=����x#*D;p��l�{
�WLA��V<��N<vo\9*�������n'���m�j\)�D3�-�J�r�0fLu�C�euWM	q�D�B��Îe���t�M⾐s ���()B��_Ʌ�����`��u�~@v�p�F�8?���	����F��Jl��u_������ϻ�骓X�t�
7�M�iYb�?������a�kϠq2��$D�!��� �}�dWn���t���7�Ѩ�y����E;�y��EeK�"F����|&�N��'�2��0C��fY��B �P�����X�����jX��wtz�.8�砟���Q�6%(C�H�F�M��1"�ŅP����80��4|5�-N�00��5�v4�W�Zj+|�� ��}���Z�g������ı"	~���@$(��{�(^{�-Z��ؑ�����K$���3d�cd����6#����i��倡/<��7CF|��X4m�Þ�A�xb�WP�D���O�6h|+��W(�p�՗�⦚@�^�#�H��CŊNp�
�'�%�x�ջ�y/��;+� �ŏ����V��	�!W�A�D'>x;����a�����-&VI�S[%v��b�b6� �,�.aE>Kgc�,c��A�_��o��8���K8��,�O���CX>�N����1	I�����������l�j���д��7ǰৃ��*�X �6IE���x�#��>s/�+�jg���شu?gb�,x�n��q���
bB-���D�1��Ag|�u:f~���6�˝+����ps�
��A��1�B-L|�l�y��	��#F.D�\�A0�������hy0x�R��p�Y�:��l$�|���{�ɗ�h�AԬV	s�ނ�Na��D�D���[�)(�e�II�X�p�ˋ�T�I1�s�B��m��,LO1�m��Wy$���ހ�cּťf���.��d�h3�q�DMg�J��N3���B�=���"��Cg� Uv�A��q/݅� P�$8�X0a�/ظ�(��ZX+�Ч���vR�ɦ)�/4��y*w��O��~���20k�T����6��H�y�� � o���G>ޜ�5�5o��g�`��?�L;ܼNA�uQ�tޙ�֦y`�;�Ψ��(;_~�	�v�+>��g�ʨ�Q5	��\���Y	7��wc�̧���6��\����~�;mʅu�GdN!r
��*�����e��ja�;�Κ9�*�"�f{
��L�OC�|����g��w�|sؽW̕�%�f�hz3�o�f�"��Ҋ��:Q�H�Xr)�E�X>�$��S�!��u��T0aP#��t?��v5���3a�a`�K�UD�_�hs��5���H
��,�ۇD!���y<=�g�~9�.�ۛ��E���' �Ն3g2�v2�>�Ʒ7��N���Ե��ޕ+�G�
���M7e5���Mj.?mZ4Ľw�@�x�D�ikp #��tB�$�g��V��^��
�r����[��Q/^���I���������Q
�x���P<���STMoVә݁��~����D3;M	>���:� D]a=G��L�&����o�r���`~<K���-�|7Hc�L,�W�k�`�#
���A�M��qmp����o`�������8�)>\r�mގ�BZ�����������-G��*2����>�t�����0���r.�!���kÞ��{�v�>��V�t��We@�B�T�F]�D�֩�W���7�bO����+p}���5�����2�(X�~�"�Џ�n����S�u��Wf���=��7��}�3�Z�U��)D�X�%����M�xuc}�? ��o��>�qp:y���)�JYZ".�j�X�~0�μb�ӹ0Av<�6Xc�S<9�V��בD=��P8}ʨ{��z���c�r%��2��f{F��Q ��Ϻ�ؘ�O���a����1��� ��q[��i��?=�����dx�{�oEy��>�Wۍ��  �D�5zMrb,�'1���!��bb,`T��(��Q��J�}o�m�5�f����f1�lr���{��/?vYk��{�Sښp��Ǡ[W��ѯ��աP�H$��=PC���\`!�t�2�b̩G��6�+_��uM�z퉨��z�ch�I4�X��-z�ի���sg��e�������b��f�Y�q����n}7�ѬőN7�[}5�LNf���d���٘�����3zcƓ�1��9��H�����8�'&�p�;��"�}���w���,��s���و�yD��lT�
 Huv
A�qw$m��{(dp��mb�)�V+J���9l���g&�܁����RVo�ō��"]KS`����pbpCj�h0ۖ��~�ukC\pǟ���Ǟ�\}����u���"�t���ڽ�\8�	�>�U$�	���������c�1�� �M�vܾ��Y�_>�M���>�L��� ᷼��2�2��ѳ��Z�i�/�-¡������'~�W��k�
خ:����%���X�`Z�w�Ǳ���}/���]�Љ�s����Of����������|�5�/�L;�j�����`�7i���f�8D�)�k7��+�}�1*bs�Vj>%ĢP��#S��'	XKo��afM���ч�{�ɟ�_�^�#h߷��A���CJqF1�Je��(�Zгk0ᢃ�ry�_�0m����G�\����S��bA��w$v����N39�j��f7`�I����ѵ�Ud}`}+�����ݹ˰^�AU2�[���p�	?�N;*��������}
�]�~;����{	���mo����c�	;�Gf�/��G�����L�:��ޛ�O��v��S͆�p�ч��ú�*4n ���	��fu7�;ءg~}t?<��\|�,#�	a9/�	�.�궫�}#\A�`���B�sS�E[�& �H���JIP�m���`l�v߸M�z��^��-%
$j-�R~{#�����:#W���,�N99�M^s��$�V~��c�S�(����Ba�n9�B!��]%����L��B��j�Վ�ֶFxe6+� ��Ч_����-L�d��e8��ݽ+��V��oB}C'�c	��[��Z�e�䠐P��A�J�V�mCn�h�&���_��J����:\e��",听�C{فG�	�w,Q PmG��E���A��p��X"H��E#z�J ҜiT���d���ɷ�:��ߝ��wf���mM��H��ٔ�*�3E��@�z/�4�vL�ep#�74��H�P�\�^��"րnZ(�J�c����h!�%O����8�b	�W���V�%�h��ajUx�e�ښb���2m>���t3&���Dܹҏ���X�d;��x9�c&JtR��(����F�YJK�P�G:��lG��!���x�$�fR�|�ݲ���	��	����Qj�p����'��L-E�dmR�$U�n��1���1&�ҁ���>���9�����y�d��$-�N�+'acȴt��dWA�-�mn����
3���G6�!�Ƅ��#l(�uUӰ'ס�x��v�|*|�Y�ܶQ�J�S�6�@��]O�4x��\�\l���<�I�7��䁍�z�dP`K��""�<Kn<�<bF�ؒ���U:���(�]L��T*�#�E�"�� �]S^�	�� �u<(� 33e�Q*�?C�1Q�d[M�s���!�������7�CH~��e"��7آ	-����W�oƶI�-��!��u��x>�)�f����6TgMԷ�	9I�o���p=f� It���/�1��K�G�[3\yR��!�nh0��O~��9��Z䒭X,J��m0����.�E�%�տ����!,g�f��R�@��-@gG�qHt���'�uHPY'��Qd�P���E�;���|^f�cJj%�M��tb��N�,��QN�^�ȖCՂF�1�kW���c|��h�j�(R���K%��ǶL�t״b(]xAI���'���Ϫ��L�$�.�\oe1Z�IV@Wz�P��u�✘|�i(���h+�$C9�	![y��W��1C�AQX~Y�wT[�ZaHU�DL�e'��t����d�"D@6>Qi$�9���Ǫ7�D2[�Q"��V"�A�U2��䁂��#V����y
�<	�0p��3�U0c�eP	 ��ј�R!/*ER\:@�'˂K{�h+�u������|f&�|ɖk�)�>�_C/������!���	S�±SR"��v)'�1W�c�O&�-����8�����)�D&f_6�B�3����(���#H�g\1�q;�4e4��T !z\�.ȶ��ݾ��:L�$�/R�N�W*"��(�����tH\���ֶP��4D�e��W��u(�T��ĉ%%��R �%��c��]Au�A"��b�E�ku�ĥ
ZK�����\}+�C$j�F�at ;Y�t��/���FC�����nG�ן�~���Q�Z�+��. ��z b��5;���Ү*>�~A�V]?�=IU1�s\d�H�e���e�2���B�g�@	����6����L��;�z�=�tx������.���%[ذu9rm+�Y�����(R=?��J�Z���1��}7�2Pg�%C�l����X��2�f�`��T��mҷ%D�+�E���kuEu׾(���ld��I	�-�L��.A�V؊��M5��{������P0�P�g����ڜ9Њ�Q��,�
ꊆ(�_`�`����m��&��D��bB����R���>\h�*l��P�{ �e�%@Ls��rff��/�EˬH���ƀ(N�DgY�`x����]8=�����Ku�G�9W�e���p��b+��J����1P΋X�D��=����s�bS��?O���@1�������2�����S��/ zFv7`w�@c����z����8��?�4�1�W���G	�s�E�O!Ձ���$Y��I���f�E!�p��Opc���Q(�b�LԘEH%9J��1c|zǿ!cXAU�&|6����cp��=�d��|�vL1�\W���$V�g1v�8�<���?�F���ܷ�P��<�|�ƣ�g�8%�(f9єU|S8�=ޞw��{s�ԋ�q�Y�b]P���!08����8:mh�x���q�Ǡ�*�|�m%S���W��e#!�SO?�O�n�.GCeyƓp핑r$�"��,v����G�+�����{�$z=pᖋ0l���'^�����Q�E�Q��fɑ\��������gb�������
��I���S%-�G#k�����%M�v�c����T�� 4���cף)B�JIԇ-�=����5�*%��h-�u�E�`�Iا�g���b��y��ȼ�I���/�N��A��P�네3�����������1��?�� jw)�(k��m��%�$^�KL��"{��)�,��z��~�~V�}z9M8﷿��0bP��,�T�B�d&�1��'��7-���+����Z��.٤�N/�ӗ�Ð�&��ݱ�9��C�84NwI �4�\WP�0�x�Y��4���9��i>0��5u�$^Z>k^y��]/L�
�U�]���CA���j|2n�n*���.��H����2��C�ƽU��i�!l&#s��K�<ߚ���s}y5޻uι�D�kI��ܒ~ԨL813m�/�!�<�*�=a,�>��Df��������ܗ����0��?������JA554���o�|�<��d:������mH����t
۰���7��O��� �BG��XX��bP���G���K��㗗b}P'��m��˷�������0(���c����������%'�(=�׏���=�qH$�N��P4ѫ�����������a�%�����A��(��TU>�|>n��A�7�����#ű)]�(橮$��-iW?�cx��ؕlm`P���	W��O�A�v�
[�8�}��b��n��n�N=�bl�a���@ul��ٝ��r3
_��E3�Ľ���sr�^!�G�w��C�������ć^��LC#:��'�&�Ð�7�?V̺=�\z�)(�R�G�l��lT��-<��ۘ��~z�zW�%�a(PL��b�[�`P|.<�h��,J�{��x(�B�(�D�������c���E:H�d�����!j�,r�����'�����Y٥2�i$( k)�Y5�v��.ĵ�c�K�Z�f��y��F�
�CK2�nz��Ç.���}+F��U�o0{�8�̟���n�R��J0d�� _,�w#��N'�n�]���/���o=����.����U`�&&
ӌ�+���G�c�3��Yw�I�8�F2։K`�Κ�[�Əu�O9^�����nR�������k�t�p	��C��rXF������=�]��8�!Α��L�GG��G���'I\z����W%��Yh�(0�Y�	nM�An��X��$<0c<�0#T���^�v��̆i��}�?����h:�esVS��9ͷ�C7<t���;:[#���训�[�/A�6zVs���8��#��T�$�d\�m��9+����a��[�&8̒�@�'�d��g�c�돠W�ZQ���O����a���L�T��M�7�1�tkD��*�0c4|���h��%���E�n�-�uM����$%��A����v'��Xl(שVT�(߅��]w1���W����@)��g9P�!+.�Xt]l4�6]    IDATZ�G���=�d������	�*0���#��N��$!8w�]" 0��eőI�֬�2����"�r�g¢=�f��Q��#2�n�|�@���N�2��倷��ӈ8GC9"���'���7ջ��(������>���� �44��$c0�G�Mōl��z�����J�1����)��7�OF�{��K�
�*oL�����
)��j���������(��B�́[���/_�抗p����e�2��t�n�$�NSs
�W�ÂFk��߯G"�Q���-�d`�m������Nئ��BlM 5�RZ=p�$�����Y�A܇l� �=�Jl. %��g?W*r���#2Sƍ�2�ok�:�RcL��Y
������P�{u�D�^�\@��2u���y��w�ᱏW*;�$qL�����}/B�d5�$���u]��P�6,}{Z?z��6(�]`(�;Ճ7�1���h��Q�Ff���Z�c�;c'�K��!�٪(d���1[pc�����o���6�S.C[�V�y`�-�-x������
Ze�*�@^�� =��ɮ��kZp�3��ЩhM��zEށ�HW<X�>[S�B2��!c�K�A�o��Eӊ�� �E�/���t=n4�|�|5�C]�@mЪ2�_���xE�>c�I`�.�V/����tc`p���uT��X��T9JPhS�+Jn3d�o��p�a�?���Z�h�Dƽ���Z�a��b��|�8��\��v��.r#�IUk�������C�þ�C�슂�XJ,�J�+X��x��?�����f�!��F�k�1|�]x��T��pK�:�)_)V7k�.�:̾��ck����G�Qbjō�sN$%}tbYj/O�	�l��$1� �Wc���W��lW[T����Ӓ1����(ql��0m�?̞�k�#hһ�d�Na�Д��1mt�rX��$���� �m�K=u7A�T`��AWs�C���c$0Ȱ־؆%c�k:�H��'$AL.-�?�dZ��+K�/{<����U���E8p�uh��Q�و⁰]�`nn�_��������7�U3g
�W�0�V.o���ߏ�gޏb��pEԅŪjUU��L����%Ό��_�Y�������F��hYf��c_�b�fg���eH�t |���\�X��3��KX����%RXE��'��(�U���$�%�e��֎%o݃���_6Z�o)c��<J��NR'>Da�:������-6�O={)ӤӵHʜg�{�rM��xa�R<��2|�x�h�ȋ|�rT��@������Ϸ������\ps?�M�!V�FkW�1�ҩt�d�v 9z"��Y�$,����l�J:[C8����������|�΃�=�.<� 	���M�h���!�!����K��c+qȹ�Ь�6v[��6�翈�/܊�R���U���I��r ���&��L��
C�ƣZ�ہQ)>�gq��}��{�}\\��#z*0��c�o�c�D'���*��V�]���7���'W�a�eW�)c2ǨC�
��o�\�����G�dZk$$0�����}�Ԯp�}*cc`�(��O�1�&|8�5����'��Y`l�^!v��o��Q�Q}��c�;ӱK�s?y�L.��SGh%0���3�%0z���=�Dʄ�oC2F�(QNӢ�-���}����r~�!d�v���^�"5A��*��%�����*cl)0��І%o�������of=�]b���S��S��.���&Vn���-#�g�X���^�μ�F�ZLىs���$;�%,z�VL����ƈ�π�-�-����vu#.���{xc`���f<�X\	.�v�0|[`�;���E�?��x��r�hp���ܩ������Ģj�x�k<�\#�=��#�(Q`]���7����W�A�ƨ����/��ƚ��(r�ChO@��*���/+̐�f�(08����qS���?[|n���]"-�h�!����(����ͬ�%1眰?b�n�$ ���R���T��*O����ԂCϾ{��0�!���ƌq����I`DXN����5\|�r�	�"��� �U����c����jծ�WG��q�TsW���x�Q�nǏA͎Rn]�Ս6!d%����G��g����sc�*����yMܮFʽ�I4�����7�`���C���f��l\.�L8 �0w>�~9�A'AZ�vՐ�j�YƂ����g�boh��"x��U5�㢫H�.k�x���x��=�FlM��Kl�.]I-T`,~~n��<���;�!s	�j�F����hn*���f [����*��H��H�[�0�%wt0clu`���u˥���׮��
�D�@i���Φ
�@����	c�;��D��Q&G�z�Da���������̀p8�D���� �L����P���^8`��X��;aœ�������q�0�E����J5��X*:)�X(�}�tv��H�]a�`�� +�8u�,���ͺ(m��nQ�{8	"A��ϙ[9Qt=��8=!:�$o3؜@C����YX����(T f��m:x=��*��C�`uƐKF��[��U����&�Lc����P���1<�!���|�yԖV��)�����Ñ��Ќ�4�0D�����}�DJ1�`�̳Ǣ��Q��"<V�q��d>���.���OM��i7�*ge�,�]�����cq���LL������bu��0�sՈ�4b�<"�6`��5}�+Ǝ���%]�D%���2�MA4���<�����Ϯ�t�d�Ő/;���JҘ���(��Pn�n[���^@X���iZ�(�C�z'`�ð���G:��lR�}�cA�xi���c���&�8�%J|��.Ǽ�1X�eW$,�FW�>�N�]	Q�X_P,(����C����FW����/��'���iׇ�,S����1�D!���:�3�^��'\���{��ɹ,&wT�R�x+��WON���7���&Q�m|�Es������[31m�+8l��X�s���+�	��t�f��wr�?��7ހ�����7��6��$P٘��s�˜����[�5�����<�q�bէ/!\�
���2.��8
W[e��{ �F��W?���b�翇"���)nw	��׌`�{�������"�N����^�!���������и�<���06X=�JMXW�*2��i���d�E��[�]%����s-~w���>��0�O�N�-Sp��G^	?DU���`�IW��;�:���g���!��ފ���wb��7
�U��h2P	7��ƛo���z��=��t����Y6���d:�����B��R����:�nM�|Y��1L�Y��4��^��F�b�������ki4��+�_<�i׏j �°�
�Vf@9ЌLC�$�>�&^��{��9(�c�-M��@��_��z�VL��F$��rW"Z>r"I�$�S@��͝����C.{��9��_!��5�%�a�n(.���YcL��#r�[�J�x��
sf܌���$O'1���Җ��%��ō 邇sG^��']��n0�<i�-�Z�Q����]�}�nL�~���hW�5*�c���)+���x=��>���]ap�	��j��Q�7���h]��p�h$l�|^p����@��`Oa"``<�>X����^�f�q�\� �]#��x���9o�<�\{�Ŝ�tX1d�98���� �g������
{��TC�E�s%�"��E�1wL�Ն+�!&��`��D}J+-`���q��ǰ��I�$���hZ�0�Wծ�����gv�͗oY�sk�:�NF>��z��ȁ8���D�F7
��ȵ-�����$�<�Jl�eH���+��LS.\��
2(�x�w30�c��K��z��2�$*q�iZxc�'x�Y8�;�����?d��P����P���/x7����F�����`ծ�M�l���䳘��Z�s��h	����h��^��z��(~����r�6�P"�1���J98Ҷ�¾��ԛxc���q6�<e+!�L�N��O�[��>:�M�*��R�n�w����Z���/>����u�DdR��Xr�P�&�3c`H�U��]I4��Q�52��׺M��;��z�B�{��r�>��
�F�1�k��/F����(��7����OF;r+>��Oލߏ�f9#P>���� 
1z=��{}�'��9�;���e��� �8t��zvγhZ�.��L� �`(-�1p�LN�3�^���Vf1��ñ���G$��47���_�	w�L\s���͍�M��x2&�~>��GJ#q'	����xk~��rZ�*xvJ�	nbƬ
3pW���L���nAJ��&��h\��|���O>��w=�C/���ZvJ
Ve[�D�,,�EeC��H|�ٻƏ�ѹg������?P�ٚ� ��m�g�4/�P��\�7��*��h�����w�����"����5��kHy�W~��OL�,@9A�0�s�����
�ͦt�{�~9�5ZY���PS�;�e�9����y�)�
�z\�i*쳍>W��ό������3�E�������O��Âw_D~�Ӏ������Y#�+�wJ>k�w���Yhu�(�D��`��D�5_�GJ,>�AQ�d�.�]�l�M�����7!��A�>?$mG���䐋-�V���W�(��_�PfI1�*1']5"�Q �ݪ�!w�SP�����p�6X�Cw�$C+�JǮD�v��m��I&�Id�:x�S#=O�O��LCa���3(�����Př:��� $7��L:-w�'��������H��ڡ��dh&��� �K�X�{ ���q� cA�A��,�X��6Ӣ��+߈r�(礫���RS���&
�r��%��V�u������T8��3�>F�Av%�]ݚ�PMlK��s\�E�vQq��"G4?�c��Z93%�����dh�	�D:�t!��%�>DBHɂ��Z
�h,�(g����F�r�f4Zbmn�'{J\��4	�ȅ��
�h9+%�9&��X�j�S�G�\D�C�D�R�VY��5���j�*�[�(MPC�5��,^U1�4�*���G�Q��5=JF��O��K���HoDv����F����N�����KYT)Zn��ۡ��QZ���O��dq�)T�@���``�W�GR�\`ZaF�!'KD2�7�!��vI�óU<\I�*?4:-Ẁ%EYC��5��*Spefǉ!� �d
�� s��nW���Vv&JF��7C��L��>8�si���wM�2�4آ����
��+�X4VG&�Id�DEHyK��B_�B�b�A�N�&|<���qc�lή�a�8N��LJ�GE֖�O8J∁$fp*�q��񆋰�����	�;(F�h����E�1A?�5��Qe&U�(?CYw30x+6mJ���r+��H9Ϡ���d��qE��d@�x�"'�x�����H�Ӕh
	?�A�h�G?V>,q���SX�>W0��uTΚ�<�"j���=l�"J1�;"Pi��cgS`��K��e�q�O�9�w����羇r��^�p���E���+�n��7F��se,���QN�܍��<�B�r� ଟ�H\�g��cD�YX���� �y3U`��T�/t��&�b�RA+�e�j����<���Zo���yLX�|<.D[e�d�<�|���`�̈M�q�������J�F�|VTT�#Z���f��k,�~����U�%�kb���_��F�0�Y�D�v'�:Jd���?0$��jW���RW��M�'ʶ|���QGwm'���L))FUᤊS>J�J�C9�#�J��O�T]��U}Q+N��h��Ŧ��V���C*GG�1(���a�5��H��V��,<�� r��p�$yE�"_�~��<�f/Z�c_�1R	�cS��UQ-���QD}~n����/T楊�P��7�j5_��m�*>͍��%0�]��0o�|*K�
kL.Nt!7��Q�D\L�F��H-��,�<~ʏ����0��i���>E�x��,R�Qe����Ճ�o��0��]P*�D��v�v�8:�虁�T&=<�:\I&(}�YI%}Nf
�xx|H���[&��F+1:�YC*�Q�I�-�3k ��{��M���T���Mq7EƔ��*G�a�{D�I�ԋ�Ht�5�>�L��2~�k�i�fy���_���$z� Fda%$ y��gy�� WD@9R"־ �&�|�����B.x�RE���UlO�K��At�J9e>i��������.���{�*y�6�n\Ή�w���@��ZW܊����}��V�P}$�I^f&Փ�5��B6�Fbv$�������fS�j,�U sr��ḷ@�����"e�����ˢS�g�L�U�*���Z�!hפ���x�'���o"�m�#	��ƿ���N�W7����sjE�&�6�+ ��_Ԏ�8�����eJ��w!�	Ӷ�泈9Ԩ����F����rY%���!G��g.<7�H>�eU��p�u���:M��d�Q����S�CPwӎǐ)����e����ԓĖ��\����J�@��N"��Fw�جZc��0�(����%�^�Ϩے���Q�]�Q�ߩ ��3T'�^�����p��ZLJ�D�+����~��ˎ� Gn���:z	E������)�;��<0�4"����e�w��=�PB])�����/�p�У�gY	����ؘ+�q��P#E'���E*���2��)����Z?�[1�G�"�T��ȕJ(���;�QA���$� vٓ��O���,��*�b�Y������ి�WZ�ddN���rQ���ř��9Q��/X�Yp��y��ٕZf������k�����W
08�|)�):P<�|T�.�&l~��e,����}�y�:t�ɟw c�$�I���r��(zE��h��PcI��>)�Y ��E8�����l�[�s#6��b>+j8��EN�"pRhn/"��H�yT[�ީ�Y�n�RI�VR���� ��D�4��"h]���!i���e_d�S19��t�o%�C=z��rU�0Ljp� �����D|U�ln� �K�А��r������m�U��j������P����t+F�(q�e��P��ކOo?==����)�30�L�q�ЋT`�G��,ʬ���վeb������m�ߦ~����5��D��jt�H��֮Z�uO�n������) Ā ��/��^�\��;��mR3p�W���� ����ߧ�~���g����? ^���m	��~:����g'���=��hhk�@=�a���3b�Ӊ��bI����{�V�dQ(f�b�����؄��
�$ߑ?W6V;���S>����IU��to|�2 �!t�<ЬYX�q�������a�n�h�s�8��-�ŷ���wJ`���<�̟�}��?�;�E\s�0�n�I4���E�[����?c82f-��.C�����᧣*��!�=����m����Ћ�AZ�F,,�����нk�,�x\P��ؒ�0��I���@�'bz�O']�a瞈���F�Ǜ@�=��6�K�n�Cp�1Hl��}GIOS����X�(ss�|ci�r�Hؾ���~�Ѯ���Yx�F^ ��TZ�ʤwk����r:.��P󞲡8V&*�]TQ�4\ɦ�N}ae�0kҘ�)��w��n!0=r���7F,Z�t���q|�.~M�&c�u� ȳk�P`�Ӱ��9��F_�Ç_�l�;��E�;�q��Q*)�5�I���_���u9\5�&0�jd���i|t�Y���PW�I::'��J���>���$h�,���]�\w�Ht��M�b�]�_b��%�c�� �Ͼ�Z5���^JY�F��m����o<�`��$������b.�,�D��ǯ�АB3*Z��T��D���Qc\v-���<�Ja��F��^����)�H _n    IDAT��r`L��5���>A2�Fw*��qѡ4�,¦�X��͘���ÆǳMv:V�p��q8�?�9�-K���`�b2�v�w�"eؖ�ōy���Sq��k��o@����[~��:]z�Tn��}�]Ӏߎ��G��t��Pk���� C@��q���SC� di�(]�����.����D�Aڬ���E~ ��5���%T�!�~�6r+���N{��������R�t)�#E���������V�r!Tn��a5_2�ć@=M�\u�����-���F����愑�S�{�g�����.�7md��Hī��K��c���q����2� N��� vqc��D2�hKl��_�p��I��9���N,��0e�p�Tr�MXo�@�܌�������.]�t3��Db�,�4g��=~<���V����N�M�G�.�jmz�5�� ��8{�x:�7(��mV'��!�r¶��J
��KRp�9|3�֭��CQ"�?g7#�P����;	�������h��uߴ�Wˍ��7����۰��u(��%> l�"��D��a��/��g��]�O?f���>i�w%��y���G]��!�!��'5�$P�*���UBn�L�|�6<x��02=A���t��l��އ�-�Ѽ�+�߹��*O)�8+U�|����a�~�$6��	��[���ᦫ���[7�+(�H��bX1\x���w��ж��b��y6n�r(���	ߧ1�����A1���+nĮ�ׯ���j�2�L8�kg"�5U(b�ϡв;>.�n���Y�W��+���X<���+�Ҏ�,�Xl��L��r���"�Y�f��?F�b�YW2l����n���-v%*0���!N�zԉ���q]"A��0���oc��ɸ��+��-]�h�h)��e�q��p���b�����c�_oÌG���#�K%MGm"�EkҸ��;p�W�X�z~>��t�t݅���C2'��o���bI�2l�����:��bָ���G��s��� ��I�z�F\�}~zܮ��uF.�e6!$��إ5�c��O!�Ҍ��OKD��h�(��j�*���\���d
���o���h��� Q�r����2w&�\�O+�O�Ƞ}��h��)�I��w�<�}��1z���.>�}��]��z�A$��q�H�W��Ϟ�.*2J���N�c<�i�c�U7��F���B�j)>Ǐ��,Kj�`�r	�(����f�q�yi�q����O#ѩKW��p���i� �sɕr��ﳏ�-�<�R�r�p��7.#���������O|�Q0z�\�rNg���'��U�6�a��#�܂���	\����Z�݋�W�[�"��ʪ��q+�cK��nį�*"�c�U�SE��V8�72Ȭ���9�c��k7|�?���I���rƘ��މFԋ�,�Ǧ�"�r�x��JM�.��#��[P�P,p���C[��ܯ��?%��r�V|��A�vqF��[HB|��$v�y$7�(|��k�uie���+kh��;}���;�K������y��CUu��Q�.�:C<��y�=���Z]_R�������wV��'̰��ȥS]����E�����%�F��j,�\"��R�������޶�����T�&E�BU�wZ��d`�H��ȭ~k�|�A�ƉM��m��Ʊ�w�	�;�1�~75r:�|������ yq�!��2c�+^X��S� ��a`O��� ����^�h@f���*rT�*�����������Wym��y�op����g��9�Y��O��M:��[�Z���E�^��lK�r
z�,��U�R䏋�����Q��i��ŕt���
�韼8W�Qo@$u����|���H�iV����nD���ĳ�&�u���{�{��3G���>L�F���y|���(~�*Pj�11��!��Ӱi_�`#��T���-�~$��L8�ݨ�Z�ԱPR���M�'��'�X��^v���d_��~������y2�R�sz��w<���*4y5HF�'ї�3c00x����g(j��J`Tgj$��Ѱٗo�P��e��E����^S�6z�S0����QQ��MT�mȯ~Ec�97#n���1��1e�#�9���O��A��ڰ+ߞ�?[U,Tn�T=j��p��1Me�
Eo�����4��=A��Wc��z�	eSs$�V,�D�5V󏲌���B�ΫG�lu�������5?G�
:g��n:��Gl
��<���D_G}؎��@������V�By?ɵvEZR�6��Q[l�eC�yM�Q;r�ȕ�����A2�����&�FJ�^Ɗ/?��a��1C̾�ܶ;o}����E�����!QX���ߏ5��EP���iM��$�@��ʲ�B*7K	H�/b�*�XL���h���h-�D�1sk+.F�d�O�	������E�1�����U�4A����@��� �_�ɒ��A�09J*�d����5��ϐ�E5�ڕT��Y9"3G*Ҳ��M7D��:rR�����_�
C��b�QGö��$r<ʨF��D�I7=���hcq��j��ȶ���ӑ�[P\�*V~�)vv�pwgO�6��Qm�]�z�?;����s�9J�%袷c��w������J�<*�Y�������Xe���:z��#�n��Q2Q��+�o}��n�6
�Ejn������=O�f��@����y�}������������<
%t��a�p���"7�j|^q�L	��M�TA��(�@(��O�Q,{����d09�Y�T�������!(;ΐ+�2}1���.j�k�Q*����]Wl?.�X+;J�Q�GU��.i�"��-���s�~�8�u�(�)�F��vu�O�쬋�v�᷋!
U��X��d4}� _Ā~c���&����6\Q`D ���S�CJUc�������lt�AfxCd���lW��d�=���D w�C��r�(�[ø@�C%�O{��Eo܄���hZ�ɺ8R5�ZĬ�̅ׯ@�ϡK���)heq-@�m��M�Wա�~�~��W."nSۣ���Ĝ�VJ���!�������wb�"a�!��]	��î��������#�=�-0: ZDj&���.��$� LG��Am*���q�b�N]�u�V!$.��G6ׂ�_D�>}Pv������epةK7؉*�3��H!�H+�ǆ�b'KvB5�g��e̱���H`�}�Ň�s�o���Q��|[`t<c���bNc�%e�+-&Qd6t��$@�Z��������%�;%�HQ�\C�i���	͙ft���U-{�L����X5R��a�q�n ǈڬض��ص=`�ꐰ���,il��2ƶ����EdbQ�J,#0���D��Cw������"��:��>GU�ӱ�f�R�.Q�9��T�����k_J<��g�y�X��ֵrĕ2^�K<U��E�L9'lE`�O�e�!g�~ʗ�2��Vc��͔9��3�	����ۑ͵�h�[�ż7���K�h\���z����~{b�;!,瑬������,�[odJ@]�t0�^��b��ڶe�'�5�K�2�$ I[� � ]�t���X`L���qC/���m5FGj��<�E�̒#@!�Ќ\a�����n@��yX7�E��i��ð��H8:���!t��HR RH��X�f-&M��Oޞ�Ԡ�ѵ��j5XղN�
U��H�k�20ȋX����-0Tq�q��NWB7���(#�s��mhA3��%�
��ڴޒ/D���}1��Y��t�2��k�����r��q7�/~Hv�vA��.Ы�Qݝ;���Ȓs
>�f%�q����e�m�gǋO.����Lő˷�n��Bz����n��/�Ev���i���'�
z�ҥO?���Ԇ6<�G2a�-�ʮ��;'ބ��yI��v�%�k֖�������+Jb�ǀ�ʐ�FB��hJH��]|n��{��� ���|#�$��!��)�cݢYh�`�;dw|��,����pvۡ�?�ڮp�	����T�
�n��?�$vؾR�:|>ov�7�7����a��G�h�@10�1������Q񹱘�B`�5~���uҜm���T|���	
�X�~B��TM
u5lw=�~�~@[#׎�{�C*Y��m/u,Y�5vݥ?�|��;�X,�;n��=�,RH�-��yTW�b��ň�vG[����T�G��i}�X-��pI�)nޕ(��p�o��]��G�F��j�ge^�Ѻ�t�3�塃1�曰]����j`��siT�m̝?��&M��rp�mwcƣO���3�V�/+ee��_�#~zjz����?�����������I`P��(|%I��%0��ķ��ಋ�������V��^�����57��Q��in��ӧ��v���HC�|�,�f.~pȁ�a���6�A���V<7���\Ĭ �����W�m(���OD��' ^������D���@qy�T���1��Vo��X�+=�G"��^3kg?���<�r	5	wO������N�z������KX��B���ؿ� �KG�/�tt,\����wO��{�~�����p��GB�h"@Ae��E������Ə>d�5ƶ��x`��:a��Cqo=V}�:���b��W��n��X2Ҿs��x��ѣWOh�rՏ��4��B/�Ìk�X�p!v8wO�S���୆�_zS&>��G�����^#��[�%���m��q����U2��p�lW��liٴ]�pj�N�
��2Bz�S���Q��aeW`��᷿����XP��a� ��q�ģ�>���	a����!�l���F�f�B��q�u�4�$R(�6(�����e0�������Ъu������U'W�1�*�@b;h ��G����[F�ő�^�Px���j-��x��G"��.>�z^��L[+�f�&���r��FM����^���g��]+�懯�	R��*�m���ǟG���#��R��8�X�r%z����M'\����Q*�D�xyc�=�|�8�8��;�A,=�T���j�AJ�	P�N����0=jpu,0�L{�ء����H��fx��<�Za/DÇW.��ϡ�����FQhCJˢ�q��S��:)GC>O��j�	�x��'0a���ڥ'�H ���͵��@{.��+W��_��]�r��N�8�l3庐�}�I{8���Q��1�[���U�db�*h�B�3�-*G�1�߄��,����,0HhA�=~��Q����S��tX����CY��y�V$�~�N8nW;�(���P%aHc���3q��Qߩ�D|�t�@L)_D"V/��_-���O�F�w�L;H.��6Z�"�l����n�8�0�Bہ%��}�H��|Z��f0����m��OP���y-?��~��D�n��$v�bl���X>���]�{o���&��ke��ʛ���?^�xʑ����#�+#��(��T��r��`���8�����s��%?@��{�K�>�8����5B�jS���QW���1���a�؏'�߱��=�=v̙#�=��(Q��{�Rr�)W�����ĳ*$�:(�tۑ^�!�~����}��-$�$f�������Zt�^��rG�������跣�a�FOk�҅M8o�i8��(��$F\5�8�~����6<�23���ZEE``���u�l�`>�;c�8�h�P�\�IA`�!R�
}]
t8�!SJ����k��_��d�r9�{W|��,\~����E}������NҶc�U��k���w�{��B���I�
� �+�b����8���p��g`]&��:����{�r,�2�vĲd,`�HuY�%��m��]��� ��A�;Օ�S`N�V\��22�Pη�q]��6-��~�4���#q���ѥ�u��#T%Y5�<�����ѩ7.9
󾚋;@�/H+L%�l:�5+��1c��1�'~]�9�H%��RH:5���h�
泂���w	�=*>�e��g�
J��t%�(a`�e��u6�'i�C�
i���
��кA)��d'����2������Q@���I��!��a��F�iL{�>���&��=࢑���/�`��v�C�PSǒ���u�n?<Zjg�M�����������V�0�-��7^|���S�}��]��N��9}�Y�2���n��V�;�'X�Q*`��X��X�L$�<J�s���;�`=�î���Ʀh-��࣏��Gg�b1�Z2�IT�m��W'au�Zlק�N6��Wd��G�.G��.��d�D	1xAA)�TT���d&"
;¹�-0��v�bJFd��� ќ��G`�f�+ۈ;&� �}V�{������4����+��@�����|Q�3J���I����,D�.�L{�k�d/��o�E�a��M��(+oڍ\0����C�S.����Y�F��\!)�%EAS�#�+m�����(���ˮ�QhDz�B俞+,> �g܃~�C!�G�U�l[;�S4��3����1삑X�p`uj��ǀ��%�h�+��U���f�N�� �[�wQ�����dE8j�P���Z�m!0�T,v�k_�Ppې).B�!Z�Y[�̪�X�����y眂�T́S�P.`;:��툧��vsXٴ�~_�nB�� x8�2y��6���n��B���6�]��١��������1Ó��2n��u*�l�9�SB*GG�U|n�+��E�L�$	�U�as�ihI�E[q9KC�n;A+���䱦1�� \C^�0{����llhX�҂�\y�qe���>���]Q�Q�Kؐ��"i��.]�"�̒XT(�f����&��VsW+�Q�v<0�+��+��E[��h:ׂl�
;�e��)Z�#,� �~|/-���6�X�0ӪtA�����F�^�D����Э��ր����iȕ��PLCגH�I��d��|^��
G��#c���Z����
�o���f�^�����@;j{ht.2�۾ȱ�c¥�L�J��mH��D��Z��8VI<泅"z��߷�[6
���7ÉU!����T���D6���DcLi&�"_-v'�B`�9�#RKӨ|�K���۽=b�+�v�7�9���T���*�"U���
�S��x"���FÅM�����~j��6�AP2���O�B�?yM�v?�Z�Aw �MP���3��110Zڰ�?�*�Q)�"��)4/5�Q)�b#�klx����;���v�hȣ{��0�N(�<z���s}t��Kp§VƲ��E��o��Q(�g�$Cp�B������9�)�U_���}�U��\}��8tQ)bP{ID��D����E# �t�b/4iV�I�����X��Ac56l�H?e�U_�����A�9ƛ���Խ�����o�D*4�����pp��;>[�s���ɬd��=�|��aL������Z'�F
��gغ�Q|��@�$p��t@�Z������lJ{�$�o�`P�l��P�l��'�B/:&��2-2��kCiᣳD[AFGb��o9`E��=����M]T��),��;u���g_���>�=EjbP���o��j-�w��0�[r�9�L�Q],#J��-����!����4GQ ���b	��B�RSW+�B8g�l�Z��ܹ3L3%FB�%~��i�02)�LR(%�wa۴ќ/���R2��:\TY6�n1��(}��%���kW�8�8���o�Ըtᴣ�H2���>y��e؈��2�I���O���~�[Q�4O��	q�h�)�+ތ�C�,������$�P�QsT�D$�P\\�pMPuȐV���S�9�����C5/�s�-�'R9��I��0ۨ553v3bR뛰z�cF,�{��vJ�7�XDb%������5���u"�I3T�E-ơ�_q�B٘���Js�ZE����AnڼA���:����P��#�!)�lK�hD
���ɩ�}!Zr    IDATj"��ޅak(� ���ס�<�v����F�c/!����7p��kP�ұr�؆�g�G�ye�<|�2��4B=�<������'� ��,4r���ي�Fi�JH��b��%>Q�{�LD��\C{��Nhs��n��NQ��X�r�[��1�\V�%���ka�E�b�'�iH�%��d9�>Ǎ^�sRB.���dV�#4��x�韢����	��nC�bT����Cc;�,�:c2�XS+!0QR��c���Ii�567H~��f�/"b���J�4j�E}�!2T����F�q��Q	A�sX�z��'��ٹ�lh��Z��nM?�yZ�?�������n���x����\0���#.|��y�`�d~��76i�1<T?ŧ�����X��3�C�V\,�Z�J�J֜�[�3W`Ř{� H�UIO*��Q�$HH��,A�����4ũe���:�*�'�YʑV���,v�s���p�5ȥ�F�q�/�7��I�T�7�ݧI�ք�π���0���Ȕ�"� �7�2!������	�u�X�3YqJl��V����6��L���s���Qc��7�q�K�2�48�V�4n��:���S�d�l}g4�}	��~�.�]:����?jX>��^z����{9�ҩ~;x�
1.�v�6c��?��g)Z�L�l;����u"���w����X��I�.Z,L�b�Bj�^��d&I�`�F�4a����Z����\1���Dah�G����D�����%�6�>�c��3М��J��[�y��4s�&��_�Za�%D��8��r�bK��bPI�Ee�C]���X�'?�&�y?�kN8@���0	��g��(|�7����'����"�����~=�{`%:����7�v�[8�2
5c�	�o��g�P<��M�بu����h�[x���h��v���J?���PY�#q	��Ɯ�%E�J�j�>:�.�.c/@"!�R��"��1�o�y�B�R��\/'�=���>�y���͘N�3����<�*lF���N���n�ZcU�2�A߃�*��GEf�al�S��]�*�`1A�B�)wV��$���/f࣠�R<j�J�ÒԆ�S��N���b��	�ϛ��	Җ
U|[�m��`������q��}kW����@mFów�m�a,}������Ѝ2RQ��#���PD�[? 6��C���,d�<����%��5��kV�԰��.�?��E�+�NW�X,�6-4=|��&T�7�ȁN��G�c�^]PW�UR��:	]�g�a�+o �Wo�U]�IYBF������Z%�#�Ym����kk��� ��л�~'��f���	�p8 υ�j���EMW��|T�5_��";�:�ݫ�nb���@�$��*���B���$��T�(8� �9���C�ք�����3�ǡ�:I��n��,�nC���}�p��*�}�uq�lT�����x֞=Ʋ?�FOX���/_&��je�Z	�pa��3"�׿�w���͞�Դ$l%��i��E�dS#���f���S���5����a�U��0(�+�S�j�ç[��>uN�t5�tG�yr�T,Zp�w��iQZ�q]rz�6�N���}6����񻅓1�4�ثtS����*\�pp�sp�)g��r��.؊p���a�O��6��w��
[����S�#�D�DAY����P-V|�(?��
 ��nI>U(�5p�����bOĤ&,�P�0$f4�]e�%+_�߆N�Vl�`%��9�׌������6WF*��>��^_�A��$�}�s\������|��vH>������4��G_~���
^	Y;�XD3D�����_nŃ�_�BQ1�f,�b���m.��q3N�trF-�������Λ-(���g����?ؐ���ޅ�_~���T���E�1o�$t�I#�Pq�D�lW����&_�#�}>r]C�����K0�dt�Tˡ��&�ob��M���N85}��Mn�Q%��|"�闔G0,9���(�K|���1ĵK�h�Q0e���p���H�n�H�͗C�*dZBHk�XT�_W�=t�Aa�:h��H�p��Ǣs]=r�2�ٯP�:�G��g�J|��5�q2v��n۰t�{6��~��.7�_w�FI�D�M3��<�a�5���g���y�����Y[��r�J�̽�;�Z4uȯ���~�hDl�H#)%Ib���ֺm��{pԴ�تף�^ċ7]��7�E����x�#]�@Oa��Y�u�w��_J�X}�E�oҵ[g��s���=�U�Kf-�~������{Ҍ��+��bpfE&q�
���5O��-[��E�D'����+Sb�J�a�e��l]���b|�{�y�'2Vb���f��H ��BQ�yL����	6��'�|ad`�����ա���oF������8h�I�_����ƍ�8��Eبգ�
�vP�-�P�|��>�w�0�Q+ՉC�t���j����믽�\v��m��-�_�1n�5J�V6l�#�"����<���n3mևu�E3^�w���.���$&�R�t���ԫ�����A���Î�xc�EXx�t��M�C]��G"�9��%8�ĳ��<
[�l�c��Z�J}��N�#<�[֭E�#� ��3��Vj��<��	�+��V��Vd�w�w�{�%C���B�t��;�e=�7�c6M�m�nwjPpT�>y���M^$t�/�~y��ym�J����GO���._��Z�f&Fa�=�ϡ�����"}�X�a�)��]T(��[p���PHw�֏V#������	pY:<^)�k60c�8|�4��BU،Wg_��s�a�n�%���d?�UDhW�҉W���磴�I�Z^�sn�=�;�*��I��N-.�6O=ѾG�!L�$�I�Q
)��X� nhH.�a�Q�t-:�_���q��:��FIr�\�l���Y�ɍ�E!��0!���L�72r�U\�-�e�����'� �����+(~�	����v���>��1q�Ͽ>n	���a����&�{mڀ��e|��p��W��K��b��YC�N�'N���hX�.�=s��8yW��-#�P�t�R;e.6k�P�f�2�GX|�4�����R�F=8n��3.�<�>���Kxe�0,�?��v�N�&�އ ]���N<��ǠĘ��(Q3�J�LA�(Sn�LW�����~��ʭ��3ɮ4R�@�XϬu\�C��r��%��]�N��Ft��sa���"%)*�3�JDۃ�?;�,�>��g�dt����m��.nC����'~8z��=�ipI�5�Z*4�4���M|�?����Q*�15���i���<��'8a�Ll�jѼ�cl�ۃ�9f(���S����G���|ڈ{ߏc'^�u��m��6�_�����W���^���0�;������(d5/�5WL��{�iS�̇�a�Rȕ"\y�:��{�-A5"�J4\y���K�xv˚�Z��m�6��P��˔�Th,,ɧ.#�$)��)ZN2"߳��+��
nYVa:*��4��_�(xe2��]jhȗ����ݭ����t|�<�]<v�e��l��۱a����c�;o�h5v'5A�YB�¯���3u�ƈ�(T�5o����/l>`nLшJ��{�V5fp������BԼ	o, h�8���
�2`UZ=z����m�[�_��f.����ZD����W�=c:|�l�PҪ����3t�غ8�Bd�
Bt*7��\4Y�$�F`š$�J4�����.��G� jvg�3�f�r'K��L��<�"�4;+�)n��?�5<RY[��v7����5,]0��=NW���������Ġ	J�^&8�q(��P���?����,� �˴�NJ $,�z
�Z�����Z^�]#5|F/������k��B��b��.e���]�^N~����2uxF
MZ�T-�ЭC嵫�5}��r�8t����G&�$qR03u��Z(�5p� �\�ݨ��ƘGY	X�|BW��=�X�rv(�L&����Z��bq���L
㲶����cIӦăI����a,�n���Jsg5��R�� mZ������%N�a���m�7������?z֥��=>x�]j�J�P)V+ ��z�$��5$Q�y�� ����N6ZaR����
�/!��?�S�%�)Z��$�/�B��n�(�l=]*
��tRI]G�L�͗$�Ϧ�'w{��1E,C,Sig�Q�Z>|*7�z��H�$ϰ�h�[BZg>	P�N�B��������\�<ߚ�;�bi�x��}$������?��vJ������l�ǃ5zv�2��)�ѫ��)��B�h3�q[�1��ѳFL�����!1�x���u�,Q�T:��H���2�ZYk0����"�mnCJ�0*+v|��\��i��Ȯg I$���d��'�?G�ȫ�	��l�0�x
(D�{.��O�0� 6o���J>�˼Df3>0���h���|�L����K��tV�	D4��PG�v�4ĄuM[��wx�7�F	�
��l�K>���x��sQSi6�dh�Y脍b+�_1dԨ����;�Y�c�d�Q�[�j��6����6�%�i2I���>X���y�]J[�P���q:L�Z����BX)n)�n�˓��SKOk���؅GZ-�/c|�|/�&O�f������\ض	�+��<���m�ek�^��h������j���吧�x�>ue��}ʿ4]YT	�21�c���'^��_٭a�}�#g��<���x�3���5�a��C0c�.��.<�n����)W@d�ҭ�}urwuch�,�q�Γ��U�R�N����=Rv_=q�K�X�R�`,'�a��
����t�e��'�g�Zm|@��fg	� =m��c4���z7�C�b��7%���6e��R0p�$��SQX�+r�R˴�|^�x��7_q☑C_ޭa����3FM���6F���-jq����<{VTF�U���&|�H*a~�'�8�e,�[&�q,��-����8F�!-��	W�Q#���"��ƀ��7QCU��)i�/�I�
x�~�s:�*oD�zH���?�c�����<��3�ﬅNT�����P��7[�<hV�
Me�����Z\��E�b����|6/[8�ї���=�#?5e�/�j�"�a�mM��r�FP�4�ӷ�C�k@�cI^ �c�ſ��������?���RS��h�x$�Lx�\ghе3IV�Q�;D�h1&bw`�=�1M=8���֎���o�m��""����@I�3'#��.�� ���vu�c1<��lGr�b� ��ѱ��p�K���!{3�2�7�+	��BI�1b��-[8��=�RQ������d_�Ca�f?����x��@����m�k�3�J�.����s *��{��VW���{�L�N	������x_>V��P֫��G��ʆeo����R񝯖������\8Z�oy����,r0�&�RA�mNUʛ	��cP��=����8�(J%��f5M1�7W���Ο{��R	1�1�'Ti�&��r8b��Cy�����,���*!P�,F�W@my^�c-�=��0�+��R�mj،��M�&O^e���a5�C��5S�'�T�?�\d�U(�K0���،�/���D)�/�����|�7^!�iIN�XLOb���n X{�� �I �A/lDgm+�����=������ҵ��0�/b�[����,�vVD�c����������{$��'ޗ�O�>Co��ϡ0m��C'�u�-�j���0���%m���w[C؆#WV��8�d�E�]dc՝�p���ثc��^� L�����T�|�t���2�F��'(c�c�<b��8z�5�g����!й�A�+&�1��b	l��3)W�򐽗�߈��F<s�L���Km���`��X����`R,�*���롇��F���;>r:�:�ރ�/�OY���%�jh1��;X�%��b���F������=��Q��������0BW��$�e�ni�q�=w"�u�W#h�{7P\>b�T4��Wk�P�� �7�6u���:�z!o�IBC҈S��\5��H|�Y�Ӵ�����0d�	�]���ų0n��8f`/^I��P�X8w>V����D�����a�3X�a�~ElT�qg�!L�@�h^�}\~��i'��0*�mhp�f[ҍ�i���7���5����a��I�֩C�W�E%��KF�P�9�N�����u���p264E�b��8b̵�W퍂Q�*$��\��R�������q��&���M!�`v�C�h3�_2cƟ�c�F�g#O���ebѼ�X��[r�bt����܇|DF�N 5���GLG�����`i���=��%܄�w��0dEqʜ'��1�&�0D��E���T�(,�3];w��^K��p���O��N���=dȉ�B	�����3�.�c���Y�����z�l�1�I�]�<ŗ5A���v�n����DegK(�d7�&�ml����7b�*���T��[��v��y�Gv%����2��l��X��s���1i���dInO���<�J����U���ѹs�j���	�K1BF{^C�R�95e��,��]�|�^(Y�`�Q��	A`�K*1-���~��8W%���zzVP����%31n�98f`_�0�"<±M,�{V�Z�89��'�{�=��c؈��}����,�P2
s���u�s(I<F�c�}}k���h�a��C	�1�4��蓙kT>���Fa�܉�Թ{�����/�a�㹫��x���t��]�u��rfM^��hJ��	�gF�d��c:"����� {Z��C�a�2�����lØ0�,;��pl�*��[�Pr�\�JA[ƞ��#>$a���
�_(�q=�8�������+���y���2rҼ?��0T��鞮sa9�,K)"������F`��ɨ��M<���ɰ)�#GUB	�4�{����O��KGHKPTL>s�O^�c/��l/�*��M�����KbY	��'&�_�0,;�\-;(���9�_<��� ��%M)��0eo���j�W�{��|.��JP��a#����ֆa��v{�6Ɗ�;y���j�a�a�^=�1T��:�1�\��2̝;]:u�K�{��#b�h�+WUɨxs��Æf�'-��/��L/A��&��$S@B$�e�QC��;��v�-ư��w� H�)2�j�~�B��w��/����$��m,�V�z'|U�=��r5f
����/��.إa�Y��QUI�p3V�qyn���C�8D��G�9b�ܧ�b��P���Y$WFd6�mF��1��l:�q:�Lnd���0��F��tT<���Y'�de�7��s�i8��d�@� �|��}L��z�8��ӽШU#G!�te�k�#LH�T�S�J8�a�T6���vu}��q'�9���L&��،��zl�3fa��q��_���EQ9�O�馛��悔ޝR(����~�1�8�7l�5t�$t?�:�z&FW*��8�!��k���RU$��p�%��vø���O9yޟ�j:�N@.��%�!�/n��gxeŵ����9EN�"L8p�Uh�7�?<�1Zݡ�^E�E�
A�AK�n��à��(,���	��&V��o8�G���(�(h\Z,�{5z�$�P���k��P�ʎ��ŋ)#QH+5ZQ�$��8�r#:�#8�6�����e@o�ۧ^PhZ��]�^�����o���JV~�μ&O�����=G �+W(��?��ngM��� ��p]�7$���{�kk�1�m���؉�L�����$� �M�8V��	�x��o��A�l����2'�B(�Co}:c�
�o�M��\����gJ��􀓿-]��⺃	�
ƺj�1QT����I�P#���![�c���H`}
�����l՛aI �Qqh�z�    IDAT���_��@�d�-\�����m~�GT���.D�Yu�Bz[��T[ �:�u��0k���|$�&���0�$�4/_4��=��v���q@�d�+`��}#ȣC*@��`��HBƜ���t��bHJevo�sۊM���Bj��mo���Dx�03Uȗ�l��I�0��I�������A'���+��Z��L�� /@п��U�CgF���/�1#�V�^!}�+P��x�3�*q�2�
~��c�^��A��Q$a��g	L��6�hv&n��}XE+�Ð�Wo"M�,�f���<�F"x��͟�,�ui�E)��ga!�D���#��,7�\��!�/�LjP�CGI))<]�O!?�0��&1 ������)gU���9�{镴r+���*A�:4M�\�҈i�g�[H�j�c|��j�ؾ��g�,����6?=!#W��Ie�FI<I��\i�q�;k�|��}��F�rAC�)� Nt�Q#Ur,ͤ��y��l��(��%7���![�fkP���?K�6�} �t�pG���2'�݌�܎������??	I�)����"�|aK�Q��G�c;!�8A�DȈ6;�b�x���R�>����+8"��{��q+v����x�$4
�z�X��uJm�6@������0ڄ�jWUR1{Ob�Z�Qw��{&�+�2d�c��I���Q.Tx���(V�� ?R	�Z�yTF�����.�X�����_p����l|4��7�#Ij�O;i�I�T1�ib�\�?5*{�X��%����0	K���(r΂iā��(�[b;3�؃%�n4.A��Z��\v�lE�m0�ۨ0���+�xbl�c(�yk��&�h_�+nq��i��#n)#����f�Ҫ%��!��̡x�=�:�L�S����Gy �V�^*���X̋k%��l�k�ZO��c=*wGMg����Crbe�!�8�I�+�Y�0i�'����sɼDȢ��Ğ�>1lz	~�xO��U��k�O�?!k���%��Da ^)`4y��z��%$w��hLP�x����7Oo�-q��J�t�+Hnl�	�I����O�ѿH-�<�J�8�����[��s���-�S~�1���l9^Ib���mx���-�ɱXFȄQ���v9ȚG쩨%ƽ?R�
���q�{'�xw�bj�4}al��"U����h|��]�֯����cH����ю骂ޫ�͆��bɆ$�'#n�8����$i����\kI�*�H������_�Ժ�3$V�5�0�¸�&�^�k8DV��	h4�c�v%�xr���Q8��p�̟a�+y�R��^J����7Y�ja:n�����!���M����r��GM�G|�$�k���oF{��u�j��Ee�-E� �zc���B0�`�Eۑ}ng�۟���M$y�� �a�?B���a�aҕ���G��� �Cl��&qd퉇��J��1q��i��ai�����~\�R�Dr8Z_�T9�G%{}�o��j �S���{�>Lؾ%�r��x�v ��tQ����j�I=%� C69 |H���sw������#_�8f2]�ױBH�[�Z�&�=.��	��!���7��"Yud���?�*�/���]hh�5�RQ8�T*\1�������D�5)��sԿT�Ί-��Q��ѹ�����i���%� Kj�4��%=^DR��� �Klb:�|���x�<I�J�h�{��H�2C��[��S1h��e�P��k@]M��7�(l�WjĖmM��J�lMg�k:	�g!�����0"�?[]]YH�]=$Uٴb⑊C}�@�Z!�X�������
ٶ}v����[�ў����D�/u3x
�z��E���!���FO�|�r��b-yF[�dL/�=���Q���lpe�r��|Ԛ6�}�W>|���V:=�b���PW��|�lY��"��s �p:����EIKAKנ�(p�>�5�@k�QM҇V}�=>�V_�ŃQ����`_��a���}G���2��˜C@0��|+�B�$S��M0��	>���J�RNO뤬-��g�B�LF#iH��뜩�ѻS5>~�oX� o�N�C�9��?2�(����T��o���<�L�|*`T��w�G�����ed����2wQ��˅�(UM���V���*��dUA	ͨ܄��%�b�P@�<�����ٴ��5�$g��)�+w�U����ln�)UwT>/G��IC�|�q���m�z
��ADb��ql�?��*-,�n8�����r�=��A/�?������Ko��OEV��hI`��#n�y�o��\���y	g�v.��0q��[���g`ejĚ*�q�h��jy�Ʉ6A�WtYHRO]��=(
�?�+Ir��*+I�e�̕�Lg�/���wa)�9�P�V���/.��'P���z�s�L�, �ƢIĮ���� r|R�U���^�f�\�V�JbFd�7�ؖN0INI*�5�%��n	�TVi#��>���/�A�{��A�^��|�����8J*���x�u��w�Mx��_��3�g�ES�F٠�ԅz�Xצ��LZh��*7��L̻U���DtԷ�[��͊m�u� s��?�.S�(f ������Yp�(e�~��$6%gUj��G�l��앴u���7Q��B�D����	�1�����q�_�~{w�
#Ij �8VUa�B|�������Kg!_u0rf�����_�� w�L�M9!ZT�_:��D���t�6���3p�����?�S@A�n
��KQ�����c��]�#�&��Il�\ ���ab������p�����썜Ü�BT,�4�� i���B"q&$ơ2 �2��HS��o~���z��z1��W�荰�֌4��`�y����t���+f.�~ρֽ?"�k�1H�Cq������q�=YjnSK�=9F�㎉X2
:v�(�x�iȌ�;���ΤMB��0k�|{��(��-A*��ܹaȅ�E<�� �����b���~�c�d�_.��tQ�	��U|�e�Ðe|�ylj`�S ��H�	�-Ǐ��)�6��}�L�N�)���mt��*aAP��(��sE�.�QS��m�]3V��!Io��~G+,�y��T-�����a�x����w�1Sh����v���6�q���׈I�~�6�N�<�mKf�W�[#5�	���J薘`q&@��isp�%W��?Mz�"\߅ǐ��������۫�����_݃O��A�=�8,�,�>R�'�$7R{a��#�SÓ�2��m�p��9_�*{�t.���vE�PVd�%�?(+��D4QRV���e;C�� j^��<��*��x!�8pX~$�y�XK�Ca�:���F��}4W<Fblʩ�u`��6������NB�q9	�j9s��@o��L-�{
���l�b��K���>�2Y�yD����qV�9���c8���Qs�D��hLt�<aq���0�fv�K�{%1U(O������б8�F�kz��;�H�J�TX�e)Q)x�,qE�<�����̒i�l�0֯�0�����.���Tʉ
�����𑳰߰���u���a���ѦPr�̾n��o?�I��� U�lI,�t���\u�m8���1�r��̮B	2��rR6B7��Q�������{�ۯ/�(�u\��\�����4�*M6��(�"Xr��u��1@fç܀��y�8l���,n�U��T�Y�HJ,)�w�Ie��ft
?�P2��0�O��&��S���)�:m[�����=�&�z�TӐ�_B �r�Ģ��S�Ю�+7�[�ᔓ���C����7Pg����&+_x���	��`l�2�T��0X	��rK�2<8����W���'7@��,�=ߓ0��_@�i��f�3[��q�R�_�#���z���[ߌ��"��Z��\K��e�Qs�Ua��a$ɧ��Y6P���Uۀ�,��C�; ]�j,E�O�!S]+B����1��_��E���F1Jn����F���Sy�Sǎ� �5-�(���i��
��f�N9Jw�c����CGLG�n����W%1�"˴z� �ӗ����!,}("�"qMv?�u��P�Jܔ�&Y�.RQE [�Im�F.q�X����<#�����G��'�1�J�T�'�妆p�;�p�1����UF\�)Ɩ7��7b��a���0�PE�43�|��!o�*��e4�������a�=PH�:@�!�_���ʫ�[�y��)�^[^v����&iZ��%�T��(Wc�3;�Aя�1چ�K�`@]�~��iP`�/5�Pq]�S�'��G�N����W�Jꪥ靌��G���[~���?���3�e���mT������d+�&&9Cd�&����ܭ�����!����o������,2��`��iZ	f���9Wi��%9��~��_�EU�e�%mB��}��?9i�Ͽªą�N����j�ap4E"�,t��`�/�䳇�ic+({�M���b�Hش8�-���dd�IL�֪z\T�4��o��������a�ᆊ[���2�ފ"�H�iőE�7	��7�9�R��V�4�?j�a�kS����14H�[p}�:d�?�'?�+������:eɾ�<IO�j�f���_�lF,�IB��k$i\k��˯��y�>�n|�Պx�n�BtO��+ K����&�G�v�fcG����X��4[�ߘ=���\�����E�2np%-��z���rو�^m}nw���� ��Ð:ݴ��`�l��>O,�	�;���I
�x��vx�U٨"_M��yղt˸[��Tǵ2���~��50�3�^�Ԑ"�Ꮠ@6�uGu8��jng��Ƕ�"Z��a��0�bzU�#+�j�P�/iKc��+��#3���=r���s�
C���l˫�D+�|H1�[�����n���Gc���W9��1�V=�u�\W�h�]��n
��P�\��X��/}�����C���Iw�!�C؄�%/��NƆ�ȑ�Q����+���!�ǿ��[����a4-[8��ї\��<�#珘4����0��Z�.�d�2����F��a������.?�/=Oe�0 �yp�G��8�`I��ۣW�mC��r�/n�Wf+��x
�?gMX��A��+�r���sD�p�:�Q&�9CSp�v��4�� �M#w����WV��/��6z���7O�Ƙ��ڭa�}����<�_�aD�ZG��-�v�����f6��o���ϱ�+`�]�d�Z&�n<�2)�^��*Q�&NB���H]���O��VǼ�Kqǯ^�ާO�'�j����/_����<M�`�(i��cH�о䳨A{0fh���?k�>z��)s~�V��4X���p^)�
�9E�����1�����ֽ{�Mm��}MҢnG��&Q�t��X
l�� ƥa8�٩m�H��6����Ŧ��Dyh��R�D=t[2���QU�s[r�{�8U�+��@��媅����A��4����C�Ƚ��%�S�*Q�A����
�����'x��Yx����l{�9=&�� �l��{k���Dmߣd���웴�iKF��n5lT�w�s(���헷�c����ᣦ̽�m�����M6V��i�BP�����;�G������o��x$wi$��ÃκL��>e���,9�⍕�t�yʓ�G���-˔�J+�����r5~�ԣ�α��� K�jx&s3�+Q	�a�Vj�$��S���;��:<Ɋ�����}�ހ��	������ݐ��M�jn���H��՚QW��,����z'5Pn�TO\�;J4��ka��n֜}���5U�W�}�7�]8]eK\�z���a�(�勧}�ҋ/X��P���#'Ϲ�-�����DÐ-3f|&4K�Ϸ��Ƨk^�|�����X��r��ϛ�a�Ð�;��Q�Tqf	�o� ���v�� Ҝ��O�W��7?^�,��5ٕ����H�u��Đ��7������rr{&I�QW/�}\���s���Ƀ$S���-�TrT���
!��(7�R�6t�>�SKf⅗�/��Z�Y��0"2*aek��{��Y3Q���C�J�b��!�S1S������\y����ڔc��0����`�.�*ӸBHè-|�ՋG���b٪�z�soCS�Y�q�z���o�3�^,au��Qml�y��t�Xh{����T,9Q��]�J���t²ZLՠ�i+:�BT����f�/�_�G�2KpP�c�	���G�1z����W	�����Z���ۊ~}���.�N��2��9��ٚ� �S�D�V�!�C3`�[ѱ�!^�g6�!��5a�|�x+np��#�$�d_�P���OB�3f���a���V���=ޤ(�O�Z��T���e"DI'B]�#��e�؈����B�Th�a���������/���� l
�����ceR�Ls�!��-"]���et��	����Q~�Y������j��: 5CH>Bq�
dGa˓W�*�/D�� �H�N�JRړ�=����3�l	2��!j�D��8�op��*�@���FM��ن?�t9�"˸(�}|��L
�|c�Ks���g�B�ϑ�.׸-�V&x��R�hO���,���2s�'+/����:�Z<�&����K��,)S��GU��l��Tl��<�F~��#�ڧd.�1NL���������SK�3���F���c8吽���"<Q�Z��
����Pf!RnqoCT�X��/gl'{ �����w����q�������1&�b(~�,��Pq~{sk
gz>JhTkE�4���V\�	��1��E� ꔃP#q��b���Y��9��Q�x��Ͽ�^�Ǥ�VL�~�b�I�<�%�����^à��*�(q���,���닆a�3q�atw6��Z&.�[�a)/�O�Ic�W_��OE��`4���g�aPK��t��R���Mq�|3�j��{y����?�+w/�/<�/���g>{�Vӱ$�y���J
 j���Kzs�҇0�y8f�upS]QD5�	�m	�!ق�y��D����Q�����fb���qD��Đ�+���(K�Ͳ8�[:硗LG���
�g  XՈ���0V��M��6b�ڒ|��ÈҒ ꑇN�:���"\5c����2�l8i�\�@ΦӢqFؘ�0sҍ8l��(���?%�Z��� �� S-g�<�n�kR+,*��N	G��1���Y��[��G���	�(R*�H�cW[����\5����W�u`ظk���?ǠS`v�m��HO�H|��4�H�����������:� Kⅻ����g��=��q�� _R6:�Ӗ
9X)�G�Dߋo��c |�D0�����	o�R��*�l�a�ݎ>���TʄdV4hiA*Q��s�+]�i���!��E��B l8���{�42Ӭ����+P�P�b>c�Sº��wPnB~u[})�z&�&��CD�Y�&X����ۯ��?�í+c���@$��ċ(�:�PP���~Ç�:��#�Uݱ>�ê� b}��x�����"nC�e��<^h80�[�����2�ǜ�c�)�O��f�N5B.NŬB4,'e���	�N���X�kx�����H��ٽa�Rs�]f���!Z�:��8�'U��y#q�vXF'�_<
�ǝ���<����OJfˠ�L!W��W56t�C�,�����[���V�|4�q�3�D&�Ze�N�@JREt�����+����2#'\��:�uA�\[��:��/���}�u\q�B`�����#N��&_�Nu�rQ���0����h��C�dJ������e�L��1p?�,�Ejy?R���pH�����G�B��C�1PV�Rg�$�D�uC�-I��-����&�Xq�CGM��`[BI��j�ֆ�	ʨ�c��1�t��8f� ��BK�p��zI���L����s�V�~��<|��}���ʴl�'$�����Q��/���c��*��	��6`�'�b���QX������_��i+���y�>�Px8�>��C���5hU��T�@L�    IDATv��/j[�|YÐ�'ӗR�ݍx�q���#���n�t��?�I�R�%�w���Y���л��KY5v�cm�|2�n��ضy�{�o�-�6@e��j��*܌�n�p�@�Iy5�F��җ�q�&���b�������y�NZ����M�v�N���d�@�i1ތ�����(5"��r���I+�a�6��W*ɺa�_
������ �,�"85]��)4�
"����YxLwiINQ�!�6�e��uQ���f���f��yU��'���
b��oy�3�j��+<�I�#�DS�uh�-ø����9y��m�I#�$�$�gV�#P��6j-]䤂����#���k:�.қ����0�ڽ��7kD��8M���1��*E�|~���.I�uN�q5���eW���Dl*�(-�2[�wcU�2�l;KXI�H�6f*��\�L鴃b!�T�VDg�b�Ȏ4K�)x�D�7 y�������G��v^A���0SҊ�����Q���l����Ɗ͒����7���8a�x��?z�Isi�aHqse�9�/]I��V/�aK�wQv}�p�TZ��n�Uf��e����7��s)�M^�@�	U+\���0ĿDj��xϗ)-x�Z�a�@x�Iƚ�����2%"|#�J�*��jh*9qY�����%�({�+.SC(�)�B"��i������^]�2T�`"���҆�D_����0�4%�,J�}��P����/H��F������E��l���\*�o\�p�=�1����Dn`+* �x%�)���[�JV��(���I-#�c�z�W-%��7�+aS�J@��@�`�l�/��YJ\���c�8�Ed�iY�XM�1����lPF�hq]�G7
�!��s�َ��[P�'�<d3�_c��-��n�3��=��T]VAɲ��	˟���YK6��G(�x��j�RN��H��*�P��(��0V���٣��{�����"�3,)����Q��R�,d�Q�U�M+Q+Hq	�j�t�|p�4t�!�����K�-���*�)T�.%���ϝ<��|��z�ghJc]QI2�(�6��&�@,+��Mtۅ��W'7�"6a�)�*'o����s�PQ����w��~.{8�c�ՠt�(OxL���*I���>��-9���B��)U򲖮g�c��0��<��6 uڮ�|�����yLɖᯠ<]�Cn %���{�*�bY����IOD*'5�J����I�9�O���I
���~�����8�I�TU�A�'��.zn����JA��Ϲ���8�5uSI>p_�]NI�ZA�c2:E���U6��A��[11q'��/:|�ra��Y�}YT���vF	;�dُ�eΐ�0�ސLSe�[�S�>�T�J�/���=��ۃ.��$TJ�"P8Q-���"5�u2�(�p]��Д˫�C�k��#�
!��Qln�ϕ8 �R���U�r�I}c)���u't��l�5!���GVg�Z:V�_DZK����;#W�s�0*
קw��`%
�+wI�It�p�M��JjE'�	p�����P��KlYS�_��JO�PjY�đ!��,�[U�7׀�AI1Ű^P�l��Q��N#�z�����qJ���W|��A�("��bI�%���dm���TTjB�Y��aC`��pR5ꁺEX��M�$E������VXB�a�{�Fs���	���<)���q_Z��Q�b�,-M��*�JY�dYF^N��ٍ�A�.��r	�Cɍ&ľ��d�#>������_B�LŇC-.�������+�oǥ� ��j���-t���lM5�%5��$��D�v)�3�BP'�7cl+�<�n I�%�r�H��������D�c!�J�c��X� D���*�8��\��ݺ�Cڑ!N�4:o�/b��*E�y(�s�i*GH�����|^Z	ZA<�DV+N�K�	�S\��+�2]�d��=w�l��x^#,ǂg����&�i��\��|N
�b���t�A)�jH-V�|G�%a��'�����Z:h��fb(���$r6+��0@���s#hl����,XF���Q���"��(A�oy���k{��C��*}S��ɤ��,&�erZ;B���6C3#)b"�M9�BH�g�34�]��r*�R2m��!� ��u�䉬�,j���؉T@6A.�T��G(����t��ư#zL�y�"�� n䢙���� �T-rVHY)��y���#��p�ɕD����p�+8_ �+�'*[�Ԭ1|��,Sl'R<;L��������\��Y(�Bx�S�\�衐;��P,Y����0ڷp�2k�!koE���L`*3-�F�F9����7���	U�#d�.̭nIT!&#���pɱ)�<ܮʺi�2Bu�٢���"���	�R)�~lp	P,�^��Z�\>&�
q����p#���b�ơ�eSY���c��)4E1�t�B�P��R7�Ur��*�&هm[s�4�L#Dѣa8r8��Ӏjzٲ���PE"�#�@���K�BB}i�E�?�&���P�&�ؕ�X�p�W��P7 ���F������&��0��'aӨ��oF��	���i�:��YzU��CN�#t���e��\C���
��ѳX�M�Ig�d��r&2`���.�ha��e갵"
�m��nظU��u���T�[���5Ǉ����a�a���(����1�����Q<�L�Z���zҠl�% a�C�ə�B�sa��<�xՖ���|��W�P(QۡNr(�����\tѣ�^H�r��l]�X[_�2����پ���|*:B���b�Qx"��͓��B�ۄ���ǡ�Bm�Z�������+��ߗ��G(4n·���y��?�U.oP3��zϬ^O�@��p��4��طe�ې��r���W=�[��;��ף�Cg�|�x�w�A��M]R.z�쁗�[����c�늌��J���{���O�0�����*ui�������L�]Y���]�RN�����s͠���c��zⵕ���ǀ��q��A��^��	��� �WF��0��1x`?4or��k�fK[K��/ۣ�ve(��1M;i��h흮�
��*�4�f��_@��Ƀ:�_o�<�V�
|��s��n�� �Y�a�]t�i�k�:|��'0�4�[?��}7\�����!���%Nxc}�B�湗�i<�*�IT�KRjVa�bȡ}1qTo��%��Qk��o�����⋿���	=�6�TzX{�!�p�/q�Q�b�y=�֫e��� �����;؝��h0P�\��ȕ!"jϬ��pr������G3�E��
Qӧ9�����{�O1�GCq�`/�=Ė���l�r˳���p���!p��/oA���e���^�V"����Si�k�1�i��3NڳRs;�:I��ت�Oվ�����}�&e"�o�ms��+n~~�%�Aˮ=/<�1~���y�yx�X��x�ݷ�ǣ�OŲe/���`�Kw����7�?��&�u�,�Q�A�.�uK03���������O���4�P�fk��z�zv��o�}�æ='?�� �&���&�C���ptg�x����p�����b՛y���ߠ��P�!ym���zbA�"M덫���s0e΋�|�m�+��߽Z��F��� ��|�࡬G��s����Q_���?���A)@�J�>[�T�!�7c��Y�}�y�hm[;@Lڃ��a�a(JQ<>����5�,7c`�z\x� �h��t�B���ۀ)�5�t0k�Op弋���>��~�Щ�߼?�w��7�ޔHےK��-f��t�s�˿�՛�j$��������]0��>�A�k?l+z�ׄ*�N�����o��Go�����ƕW��{�1v�i�h�8��#q�{bܔ���v(P��C��o���������0�(����t���Ȕ�a��`d��Kđ}�a⸓1z�C8��� �ࣿz
MZ/�4�L��'��ϋ��{��#��R���Y�w����� U�EDε�+��b���G��`����� <����۶YI���Y�ڔJ�*�GCC�p�)��ē:�򫟄�aXv=����N�|����Y+p�Q��ck�v�68���#�����^�S�d4~��!X�6��~�
�N7ԊDX���Ȱ
�n�)͍ͮ�p�1�����p�#(:�6�[ؿ�<_�z�s8x�!��I��}�r�y�x���b��0tԷ1�ʟ�SO��'�b�5� �=K����8��#pѕ�0LQ8����4�SZAHIM�oވ>=:b¨��r�
�6T&���ߏ��Fc��?}���3�����em �~7�$̜r/>3{!��yW��,Æ�!#����c4ߵ`�ɗ���n=���>r��)s�i�a(�E����I����3~	��	��Maܘ�8��G����M�*�0컇�G�,��	L��,<�Л����ix�mx`��~��V��-�p�����5�g/�OwGFKJ2͊��`�-s��T��{�`�E=1}��0;tG��ѷC��c��ᓟD���q�=qͬп�>�1���ﮧp�ȓ1lگ��O��N��u7��:[7�ǹ������a3�v_�Q;�Twdc�8� ��G@=ִ-�qż�q�-´I�`�m�����̪�Z����93��PFA�!16�r��(j�I~#�Ad�� )6�WQA�A��$�2 خb	2���9gN��f�ooa�k�y<O���o�o���U�������ˮ�h�_��폂�C���hށUs/������� ,�#P�H"Ef�^R�j��|�;��,
=4�_'�|��lF5��&^��lĶ5�u�ނYS���;_⩗_�-�]���X���֡.�桤���؉��(�ɜ1���h㞧6�t�f��D�T�7�@�9b*sp߄JQ����s���*6�F$�Y�%[8nZ��8	���7O{��è���
\��Ӟƙ��E��;`���?�d465`�X���Wo�)d���Ty�H����$R�Ԝ<�&����8��/ ��|��qr�1�:|!�pg$lb!���fa�Ⱦ��ۘ��i4
:uA}���i����w�+Y5��T���dT&$;I�q��ۋ/����w�植�N��l��]9�3z�聑����{@m��~��x�=��e/B���j�6�\$����/C	���5@���WS�:�.+M�.��^��/���kZ�9�ǅ��":�U�:�L��7���=�`~'��v���D�;�9�~֯q]���C aǝl�R�c �,����&�M�g�'�OC�)1�@N�[��_����_�� ���8n�Gu������/�@���]w\�ʝ��-@^PCYɚ��G,�h[��A�h�b������?���x�<J��F�����>5�t&o7�P,��%e"VW�ӎ;'��S�s�lM��w߆�`j9��4qF��(������a��g~->(V
�W���슛H��P:�+�Ӊ��M=I�yU�����il7"!�\t�! Yc`��j|�����'�_|�vN�]���rQTt$_�ݏ��~�Aꯨ>���d{�
�
EE��A�� %>oBN���\��t����2�G�>��O?a�?I�L�`%�����X��Zl���d�p'��D��g$-��u[�O�.֌PN������V��c��C�0���=sU)Ȑ�=��a#�#��S7�7Z�P��H.o����Ò0R-h'�nG�D
��|dH�D�3
�$d��*�����,�]e���P�ށi���g"9~�$�k�!H��$� O�Y��h���:k2�0-)�x��.|2R��P��Ɍ�K�$�3$�C�ɢHc�g/�t$`D���#�!��`�a�`F"[63�8`��z:Ú(�t>Ӏ�hJ�hױ�Ob-[��Z\͖���,�WXۢ��j@E'������I,����S�1�%f�4$�..�O� KBʰ�H�Y��:dL��.)YZ������=A�I��_h����Q$�Is�n�M���1H���a�SU0�Լ�?�d�ivj�z���_VGtU�\�J8Sj�;
�J�+����룣��b�ϝ���$��}�D"P�xV�	^�t�NӤ_J�K�=�ᙓ.1��~��č��L�#E�J�%�_P\�I�E�uN�3`mr�9V��S��G �hD�~^i�����iK�(E\�J|�t��n=��A�Fe�!�q�Rw�J1D�#{�l�4���N��7��*�ihhDT5� �GR�<$�s�1�p�Ej��bP��$b!��4!�#��ޑ���Sy�&��V~��AR��X:}!�u/DP�{���1�5����o����͒2T��Fm!��4L�:�&�i@*�+t)H1UN	�)�����P;:'Ľ��� �cW4fd�dd.���E�r���
� ���A��X�6��,�6Gy"�VEgԃ�y�Ds-l"f�izNw(�����<�"��$�!��7�0�X���Cد ������)��Mք���@���}P5���BGSFB�{o4e迉��f|��+p��/�q�o���q@�X�xŐ!��~��u���<ڣ&b>K�M�r�B�I2����&Rk�L�KuDVO%qŁx�|�D���PvҁBH�KLx�� ���[f�F�IO h5��s�t����"<j6����oݠ
�C9��~�<xD�<��A����뽨�	(��P�l&Q�y=��z�A�
�����T>�z<*)�O�r��i� �
���#1�I�>��4�KV-wׂ���]�8��/�:�;_Bp>��f`��AX����hx���EZɛ�"�[�E��ۣ- a;�G���+��I�?�I�a,���&�@��rX|:�:7㍹� f=��`n$�H�o����Ť��Fd@m��Jq�)��QKF�ʢ-�w�s/n�!�(��D�R��jT���J���Sg<�rIz󎞡��AHw�^�g#�+�e��&�q?�W�+1֔��E�7�c2��G�n�@a�
}t�/q7L����B��F����z�|�r��@��:�o*���/�Y��v�/�NG��)���v�N��=Q:�UR�%oefP�Ϡ�ڃWg�dvv�}#�-qc9�<�n��K�N���'��[�#����x��;Pc�:͊
_��M/a�ߖ��i1��j���9�����<�j�1�aĔ#��d��1�Ɣ�]�{&_rݐ���1���l�]��j�=����G
���$��AnN�H"�I�����������V�G�hE�\(�&�i�Y�G��Q����
ӟ� w���Q��4m/e�\��#�nDAf'�?8�l����+�-"F➠6W���Px�(��	;��,(�R>z?ϣ��qB5bϣ��ֲ槫Q�z)T���\2��E�m�SN��~���Dq�	�OX�z���l/�^�Ѳ`��K�J��,��~脻l�a����]���*d��i�J�Sȓh��2v�0�ټW}�{@"#�%T���$��΁T����v3)�������8��(�[[!��2��jtqvc��I�̯�'Jw[���d�Fb2J)�.��ec��� ��c8v�M�����yXWI��9zқ����j�3��l�db�Q�~�M�DW���^�}&,D����L<�����y3'^:|蠊{�%+F�������`��#���?�\�d�t�eu�[
|��1����^5���9��AWE"o4�A�:�R�T\� }�Z7�=�nԨG0��x�i @d#���$�G�N9v3
t"Z���=q`� �m��N]q^RC��G���Ǣ�	�!-�p�U���*Hd��<B�6ȨLGF;�{�il_�?P�Z��G
�b���)
t+-T=�b6�|��a1���,���<y��g�gM�lXt�ڃ��c���y�bh�����2���
6��Q����C�l��b�s  �IDATFِͪL�9̫�O����nGn��ۓ,��	c���+� �H�=�N�)G I�*�]�(���3]�`q�a�|,-C3�_a��ɀ���d .}��%�qR��ИHs
H���=��-_����j'^6��)9����<N�x�]�tw�����齿b��_Q��4���i��B$'i��k�][��̀e�^��L-DѠv�ek<}�*���0��gM��"�砆�p��qC��5���Ὕ�C�C�TB^sg��BQ������nA��5�[u/?�{��*�s=��B�"���9���$ʮ��
���l}�ށ:�I9��*�àݤ�M��J�Ŵ����x�̀�`6{�7L�������$��h2&���;����|��)9���^,A�S����a����"D�8��]�]/-㬈��4HE5��KW�b[&��(�q�5�����7,F��6Iw1-D[�.?Ʒ�h�y3�\6|h�k���ax4C%Z1u�N��o.it�g Ό�ͯ�n�}�Y�����N3f݋�Y��F���rc3�=J:����W;!)繴��+ܹ P�u\�#�k�l��x�-�U��l�d�c&��/N�	���-U������/�~�0.����EF��`(٘���<��l1F.ZP��*�~���HN��^��=�P(���pn��FL�2ŕ�d J�:i�#�X2$��ګ�������ߑ���c<�h�ء����m��
�8�:/t��n�+��v`�Q��g��(<:T����.��nhsH'���Q7s f_�d��^툤�+��jyj͕�o����i �đkVc��[������N�8}N;����"5�n��TTn�r5MX����@���c�:�^AM̮�0���[B�(Ix�����a5p�̌�2p����ɇ����ݜ60��1"���.��	}&>�_� 4��<]�	��e�fN���磋W�:����b��9=e�m�l�@P���IL����"���M�~�Hv�p�6�{/��LI�SX�2"8��<u��q��Q鈔,x@|^̊~���M��l�#Ϩ��{ou=F���ɓ�3�N�͚�A�f�uL��fl۾�5�L�.���aPZ*�ἴA���D�{A���%a�?�]lM�㟞t��#77Eg���`��񮖊�j��c,A��H7@���U~ �.�X0{��MW�Y	Sr�H��/	������p����QQ0i h��a�z�(N����F����E^$��:{i�h���PF�낳�ގ�0Zȭ�}o*g*��pD~b�a4�Q��>2�� US1f�H�:�'�3ҀM�O�6_T��j!
.��ǟ���m��6E�Dɉ����.�,�� d�a���M��B�F����9�AD�~�-��il�1��[�j��`��`*]�{�c�����h�oo�2��0�g�E-p-\�l��3�5�Ԡ��y>x��H}�(��"���3j����>�OйK�)��2"]ݼ;V- �Q��������Da~G��I9��Dݣ��Z�;�N��af����
���^����yX'��݌\���a�vL�q��ĉpꩽВLs5����4m**+w����^� �/��O�+uk!��%�'�*hH��->Z�J1�~�<����0��н�C��8�&��Q݀&L� �|u���LZ�G	���[ܶT�@G��3'�f��A�������1d���:f1��B� �"[%4�jc�H)�$2v�8���EB��x�ILA�C��+��o+�[#���m��~��ܾ��& J�R!?JXr����Q� f��#�[�`��k`�<ͮ�1����(YM�:��D�8F7�pN<�R���ɓ��˯��Ћ!��oJP���#��ʫ�z�5�����a!�ɼ~��_���|���WCs��~����׎'ۉ�1na܈�P�[���,��g�{�Z$-���j*�-�د�x`L˼{n�p��?���hђ��f�;u�b�!�!���t�N.�D��# 9̚Gmwj_s���W��p4��+��ހʏ6��:���D�@e�4f�1y9y��Q	9e��~�.|qT.k@�N�f4�"X�|����KɃ�^��8��g0:-��[K�si�L#�"��O�N�{�Yl7�<���?�v�r�(:�/�\�L�EMTQy���� 4�]i�(�L7 d7a���hx�9 ���W��W%̝>EyH;Ҏ��Ҙ~�T&���A��:f�+��˹/��5r'�����W��X��RR!`G�<<��~#�^u`������J��=��腨��9�XA�H�
zE	zBUO:k�<%w)PGn���72�US'����4�15ۑ�݁�_�q�m��|�C3|Mq�hV0�ɷ�)
����t?�$�I��a6\qxyi���T�aI�B��V-��ћ�h�4�4An�`����[;���)��ၥϠNꈌ�"��1m���w�*h+A8�#�bQ<INQ^�c#�qXB��d�64�4+�;*�D�ބ���F��iX�j�<,{�%Ȏ���g\
�[�~hQ0����b�i�6\�+y^nⲼ7Q-Ւa$�Ϟ��`����2��G��^�Z�0�����|��xR\�	�G�ܗ�Ӄ!"[p�A@��Y�rXݝ���P�8|�ǥ�uC'gBH!c+h��o6�l,[� �a�*�Ĕ�� �i*�*n��%ua�rFES�=̀^�j��'�x��_��_DpT ���3о+V��5��Ѣ��&+H�M�ׂ|}2�Z�Ȫ���b�7��N�L`!��Q��Lq�T�z9?B�j�?%cd$ah��Fg��h't҅�#�|4�R�\�LT��V��X[>�c�wЁ�K�K���Xt�臱G��L9��vQ�d��K`[����e9�V�!PR:쾴9DWd��Aq�����?V����n�nD�҆�X�h�Y_��Dn�%aD�C�0!�e'Y��[{o�%u!yo��\U�M#�To���A�b@�؃�����SKӬp"�k>m�6�H4�aPe�1�d�Z-n|�``�;:Fż,W��`��~��A<]�%�"�AH#nA�@?Y�Z\�S]�j` !��Y�7+chrr��Tj����ԓ|?���N����?��X0s�Q\��ɒ�	w,9cԃ�E���Jf�u=�bN�Ĭޔ�w��kx�"3/$��QUQ�1B�0�ڨ'��[m����%�B�ӄ��BS�x+�Ӊ̎��6��@wJ{Ncm�Hg�P뷇���!��OT@ɿ��,�X��HT�z��Ԃ�0�p� �C���1lu�Y��LC#V<j���%X��� �hT�1�n��qPA&4oBG�_��'<'�nu�j�n-8©F�6�R��:� w�V����P�v2L�B�Qj��Ϸ�4�F��ϙ���4�=;p�����9u����kR:J�!i�� ��y4�ď3� VR&W+��(7\)
⤢a^����
�=�Xa�@�"�m���q��հ:�Emb�ԋ!��R���0�.tq!�(�%�����ꋄ�th�@q^�$��MBK7C�P�/�+��?2a�
2@�.�uT2E�)��OZ�:�G"�h���O�.���,���	K��Q���I�Ȯ�߲A��NG�zo;��G#)E����� 	��j$b����"Ø;鬃�9�[�������s���!%^|"��>Z+�)�oA�����`0h�T�����+����l"S[����'�ev!OR��R��v��]ð�f���ԗ�!g�2�K܂�[�̟H[lK��k$���'霐�[Nz�.2qR'N��ĔBT|^�]Ng؁�0b��]�k��\��Y��(��@1�"�3�9�KA"���Y|>������F{�Ჟ+��ԃ�S,_>vJ�x���P{ �(6���H6��Ȥ{&�Q������;MX���g�|����[{�o�1�_�X��7�|���	r�׎)���G]R�GG���������X��"��@�K%=�MkIЬ"j
����}I�p$��=)}�v�|��7D��,�a����baL�����a���� E)����4�:+�I{����"n���g�Qk	�.�a�U7p�K�C�Ik�R6E�����D�d}��m���]����6h��io�)���AȖ�%�������:́h�[<��j�	[1�8���G�~�u��r@Ø����aCG�_���Upu�!�^7���&:>F@yT�8$�I���k?%@p�t���J��>���fh9[�E'� ��Uu8���p��I��Y��ɓ1��
�Ket�# �����1����Ҙ�S{��h����ѓ����θ��*B���+���D�{\�s��Һ�b^��E�Y* V�<cέR�<��dd,q9�I�ǘ���縮Q��������m����_��;������>x���_NsD�ḧhɧ��>��J�O<x�Fh��l����8���{�Et]W>�l�d�Q'��*�5ɤ��q'�0�w�ޱj��W�8�T��'a�R��;/���^�2�(��<�k�C���IP��C��q��a���85�����"[��������K;��Uv��=���Ϸ���_A��Y�耴�-��{03���8tȈl\�ڗ�;�zϞ�[2FWJ�e+u��訩�X��X��c��9cq�#Ѐt0(4�dI����:��a�u�i�C���2i=S>hH������믽�s�����G��T�u��*6�ߺh�/��gg4�j'�B�#� ʝ2�ʁ3���am�/���)SK��A�*�x�����������Vm��9�8�	��oWvq6֦5�/\�(RJ%�|����3h`tB��?�cٲe/�'��;w.B����ß������y��WJ?���Ej0�I_S��MCˆ����i��O<�L�/oQ�J��}���A%�Z��6������-����X���������yc����غm�i�T���%%W����c,_�ڱ�I�I#��+���?[�ֆQ^^�aƲ{R�K��۟�����ͩ�xm|e��\��ҷiVF�����]�x�0���RD�����0p������4���P<�h���'g��TTT������+��vdn�F�?��ڴƊ+��u���{6�yqq���Z�p�����k�0 �[RR�'��v��몪��2�O��hV��k+u]���a,)...�ƽ�o��*]-//�4�KZ�[%%%gfcs֭[W�u����cS4�Z�bŊe����p=�����ٸ���x�4�K[ƛ%%%����ُ���FO���n���0�b�0��������QB�eY"�YUU�@+��m�x�0�?�������o�ˆa��*�|cp�
\�	>?�F�=��ƮX��)]���c�_�|��0�m�16�������SQQ1����V�h4�+k�+W��K&���ceqq1-��s��kM�����8뮽�ھ�ؘ�k׎������0ލF�YɈܬ�]���0/..��{�O>י�yN+�������llNEE�����٭�h4zz6�v�Y]�/����=1p�@N_���˖-��,�W�b��|^66���bRee�V��v4=#k���뗴�Os0z(>��a����(�5��nݺ��n�z�g�e�UZZ���k�u]��3�@ �Ԁ?����(//�4��Z%�KJJ~��7f�ڵӪ���t�]����...�2���c�d���"]]�n��[�n��%kt]�x��?<=`��+~4�1�Y�Z峢�bzee�M�0�\��:g`nI����bN_��p�1�5M��CT���������0V��P�yXƲe˞�,����&�V����5�\��^Ɇn۴i��P(�m�T*�NYYY6�յ�a��y^E!��篺��~4�Ix¶��4z�r������|޲e˖�Y��DjL����Ҭ����� �G��~���k��u(>���X�d�R ��(�|��ʊalذa��͛gAZ:�&5�#G��e�ʲe�^�m�"�G\�OF���� V�\9'�J]o���ܹm�ϖ��e�Y�f͠>�����;��pgհa�f�0V�XQ��'I4k�����,���+'fk�o�sXy����Ζe��i�i���e��nݺm����ܹ�g�i�h��b�f�QG՘��w��A����$Ɇa4���U�=b�Z��6���Q%�H~��8�<�!ڃ�����92f,    IEND�B`�PK   ��X>6YYJ �r /   images/54ec96e0-e6c8-4747-b5e8-2cd896730fff.png�w<��?~�J*RF���	eTF"��$��l�h)[e%3[B���3"�{%�X�������y|���zԣ�����u����|^�}��UQ��`0����]�`��b0{�S�O~��z�?䶗�nP���}��~�+ڶk�����|�h'�gil�p����� �����𞕑���I8A�8s�$w�c�t��붥ȝ��	���1�,�w�[��à�+j�`���?	�����C�|��������>"*d��izDq�^4=�+��'svo�Y���Jy'�'��G�G<�C����"f�0���\K�w�c�����볃�==�[��;����'��ql[�*\�֓,�*���;c;.�%*����.��x�@^��b�%*�O��Q0�􌲺�r�7��9Ŕy���#��ƙ4k��2�ld����0�݅�sb܈~������[��-�oI���<��t��))q�8��"'_U�z
9��V�I���4�BK{1��ϓ��xVً��Q���)��g�4��4��8�g)�~�T��5�1�g�4��7�͑��{iz�a'��W�q琡�	�#U+A}ҍ������WN�.�����U>F�c�Gz�}HS�q�2��xΠ�^��E���礋0�%+AWҰ����ʊ�zoU�[9*�Ite��^9�ʯs�S�9�Is�����U�7g�e;A�g���ĕĬz8��f�l.P�R3G^~2�+���u�z��~B�5ҧ�N0��;�3�Yn��+�!��f�N�NKN�xs�xD��#�'ˊ�HU��G8��I�ׁ�r�+�'H֯��y1��J�^�Np�3���Dk�������#]��[�Ss��Y��?=�{ ��P��b�~��<��r��]���Y0�v�'``���q0P�a����n��w�m9B�x���������;z���߃����ycѤ9�D���ʰ�$�N�˭H�]$9�pͮ��+��"]3V�|ş�D�/�Ӊ<�3$xhc����J����=�\L���r�4e�x�E��N��]��)��ƍ��I����Q�f�+�����c��ns����"���cc�7+]���#���G��7o�� �S �z5x��	���?�T�d0t)�h�=�O�c���X��!�
�Rv��w��0�'l�Y\ %�z�܊�<���t�ݐ>ܻ�J�f�@�0!��_�6�
���q�fu9׼�� ��3b:r|{?�
5��e��m�g;G��0�uZJZ;��w|[�Y!iqV��V�V��gc\��L�4���,����.�k�43?����̺s�:V�1�c��{HK9QZ�[����_<��zT�{%�L,>e߿[c���	�
�Br���MN�6�#���(q�
+�H~���W;�g��x<T�}ʧ�|���T%�����/�b'���s�z�X�[�/������[��mo���&��kVX1�ߤ������7)�<C���&MH��g�oR)�kv�/��4(7֓��ګ��ir���{����Sw���A��{�=��S#���K�C۹��إ��K�W���+���=�}���{�����ߚ0ˊ�W.��g6f_��X���,{�\�p3���%~��݌5��Nkkkknm��v�Zs�rhrF��`��Ғ��.�+f�+�υ%�������}ۓi��57�&
�7�H��4�H�,�73���̱�;��k�w-�|Uw�����R�ISTk�iW�8�GXF������cgO��̲�eE!��	}J�������鼹��Y{�{Q3��,�L��_�J\��{󅗤�*g�G��~����3��Y�~������wv@�r3��.����L��+zE[�=��co�=Ó�����-���$T�����~���۬Xs����
*��?�~A^�T+|<�]��PS�q`�ǅߕ~�`V���6mt���^��Ȉ�_	�Y��^R��V��h��L�B=@��8�^�α����E��f��˭�<�N~�5J�8NK���o�{L��_�ϻ���+���R��|�mǪ}��?i#?ã.N>�5
xt_.I�z؋���;�Y��>�;�e���l>=�L�;	{Ӣ�?�Q���9� ��<��K�-����2[�SS����;�z�= ����鶵�jˣ���'y����������\�u5#�tb�K�<����S��$ö8֤�}U��8 ��-5%�+PMZ�Qr�h��ɤ8�
��C�Z�dXZ�-�1n뽒_�G��H()�n�ޘ��:�(˓��Ǐ���}���&�i_Ry�����j�\���ח��Hk9�{����D҈��:�kvvB�eg� B>��xp��q�;�P�r�@������td�U��U�hפ	�ZS	S�R�;Nw�K���˗�������� 
ҟ��ڙ��虂1��.�T�g�T#����$�{��Ba���Y��|<�݊���ݼu��Q�~�'�ʻ�I6W�c�g)&���m���/w�c9CjH�s�>�l��e�JO��P�*�����^�s�7��I$��� F��DED*GC�Y�#�.M�&�� �l��������cBo�3՚÷�-Y�����*wwi��;#!�aZ���u�[��C�)3^R�F?jO�O������F���_�{m���V�=z�2�Z��o��$��嗕mZ�,}���=ht�Jo:�aI�'����Kn3Zv �Btttֵ���{�k(s� fM�n���~&���'O��V\�s]��|,���.P��ò:%)������P�ë#����k^έU���c8��VIn�ܗ�)��5�J��,�p8�U�+�r*/�X���.m����R�-2��l�2ʧ�599ي#6���jfrX-K��]MzqI��
�c�υ����Hoϳ���*�����Ԡ5Y% Z���v�K��o�V=�����7�`��ԧ/RD��V�����*������P�8�-�x�j���99���^�Q�H���W�:�|�?����ɲ��p�D?��J)5T �Uh�����Ϙ���-�����'�����,-���W2ǷsQLN���f]g�����u�<�;��w��m�?aD��wd�&��Y��:����(�v^!D�3)211����qa�#כ>�����<�~���A��t�p�J�|�E߿��]��e�|<}2��#͎�$�K�����}���Į��	}4X��p��� �Ք�`�Y��ۣ�ۜ��ߐ,	�}J��:�d)-9=]�!����L��������W���WU!'�w�2��%����K|µY����\ˁ޸������ϥ$�|�k%h��Ͼ������V����:���$�>�9��^G��7����%���p�=m�P8���]	;g��6V�g=r���ų���+�y�{�h<o��GY�Xd� ����?D;䢥]�������Ť)o}2�U��S7tt�6�\ a�3��+׮��{Ր,��~��G^�d�����ߙ�K������<�����0�u��I��78�u���^P��Q���ˁ��StD&s�+��,=����Љ�������nb,�N_����o�p]:H�vPoX�p:k|��}���&bC/�4�J1�:L�r�q�PM%�I�g���P�Z%�`kk;��|��X����Z�d!�����5ҋ��f�8�4-��9M'�U���-ǹA���-��A���෧B��;�]&��2
�W�yS�45��7�;\~՞�- >�1���ˁ�z�ؕ��T��_� Ç��+a�o��}�Dr#�*��Õ^����{7�X	�D�������e�����',��s L-d5�Ml�w��o��7������	�}&xu��X3��iL2N���d����%�F��;!�ؔ��K����ȺcS�I�FKrV�9�����2�ý>��4��]6��mNR�n�<PV�y�F����?�bbc�JV��]eqߜo.t���")F���af�A�J�֣�Ku����u�קU4�߄N�'S��pBl�R�'���D2{%p�ڏ)�yo4x�"9���\��8�F�Q��cj*<�A��.E	A֫���
�v�t�5N��*�X+W̧;3S��h���0���G��o�̐���\�I�M����D�Y����6@��s�)
����Y�㢼Й`���f��;)�h�낂���8��9����ycw=UY�"c�;H�s���2۫�))�M��)ěծ�pG��d�{�4��uTU�����N����T{U�p���G=9�YF��=9���C\����;�mM����TC��l:���
ܥDTۺ!� �Bh.�;����e��u�yG����_�yCX9�����p�� =����IHr�H	{`���z��[f�@�����vS���||��ri�����)&A�я"���zŀx�3  B�Y�C�<T�O�tggB�vs?��A�	���|�2z@\���R�-�o�0�?Or�o�X�"&7ZZS�g�����G�?�7�r��=��q�p������� �������إ�,�<��C���d���g����6f��8�_"��%j�_���ݙgmx�������G��3L[+�b�{����W� ����<�~��}�]��C)&�rrx�ƾLw`l붑��'Jج+i���y`jz�k�M�cbV�5���{y���+^'8�2� ���G�����`��̤�M�w�O�å���XHX@�����^^{�YS��=�+c�}懫�7f*�3�<x�`��Y�ejl��م?�5l�X�y�|�K��w���̠1S��ٻ{z'~%�oo�6Q����%������1iGf�!""B��.��xd$Q�ȸ����:�_����x��"R\����C��Y�ع�������0��=殊}����}<�t��ǟ�H&(]5��|hq��#2�
�̌�yU$�b��vsTظ�:6[�Ó`��b�s#/��d(8��a<���_�NX��@�)p^�1��D��tW��Xck �m����l�5@������(l\�I���r�\nG,Ho��@��7|�{Q>p+��1�Vav1~z�'���\)��$19���B~-1��V�u,�|K��%�����z�BO.{����0Z��<MR�**�EN�f�\WW�7��	�8��1�dݴhs�~�rR�����i����M��<<�� �$!6�ؤ�v |�јD9�Z�Yb��Y8[�$�9D�k��y���$fuws�t?�H�m��I�[*�z<��U��X�QE_��(��j�ke�dj��Ϥ8磹�2�F�ʹ�
������o���ou�/9ɑ��~��0\S��*�u����G��jw����q��/MҒ�gײ�P�<Q.��[K���)����y�$Ο"_�p��8��{��G�R�P�7�E�n�B5�e%�Ϊb��iLvv6"b�E����P;O��L-Ij5l�R�rQΪ]ho��� R��iiװ�v?�-^��m:+h�=��Y�^���{�{�6����UP��
����a���G���#��
���:�ݱ�s�d*al\�02��<kkB��K�i\b%H�`��7 �7sːTϕq�F(X��[q��t����T�bԀ�.��"�:�<�~�[tt�~��*m�Ȅ��'�C�x�m�p�,+�]r��(�T��v���HD�[q�j�����M����k�N�����u�o��M>93SH���c��A�Z���.�%��g��cαo[NҸ�"��b���� ��U���������	�D��t^�s>tM:$?��\Y�|Ch0)cV��@��/�;r�/M1�W%� ��QSm����� �L��j �U��q���DC����j�|�V��N��a��0(��(,~8�$ʫǲ��<���K���Qo����D­\݃�bg!����?���tV�J��}������)�yir���ۈ��)�qq��F@�/�*s�n��dâ��E�Hh�wX�c�wgO��l���ƭ��cH��(��><�,;7����s�V��W,��,���~Aa�+67G���ѦWP
@���Ы���m{s0�lffF���[���Ç^��뭁߿�iU9-B�H>�?-X��5�tP�;� W~)�$gƮ"'[�F��V�B`gN���E��jnG �jj�ޠ=��ӸX �ȯ�}����B�I��[-g(9Q��$�a�9�Pj�b�����QXɽ��ӂ但� �5�������,�7z:K\��>@���%�$���ӈ��l�4a����V��Ȩ&��/���;�7%3��C04����.��hhm蹽g�{#�DFBt,�M@���|�r��_�@�V�JH��3��wRN6��F5���'�Zy��Aӕz�H>���>z䷏���|D2�2ܐh���?z0PK��5K���1�ͅ�R_ԩ���S
w�E��"�eeaf�g�t�&&-����{ڕww�����P�*���q�+tPC�p<6�>B�U���¯C/l�����+�/�a�QΓ)�_L�&O����D��RQ���E�!~����z�RD�A8��=۴�c�ڟpC���N�>�bx%���d��Qy�M {M!�P_)Y�cYLw��W���O�AY��A	J�:I ��IcD�h��bZp��Qd;���|�"T��)���)�[[��M�bT#%��]t .� ����t�BL�7d>�je�f=��qA�~��V����Fπ?H@�v#
1�͟;ʑ�-�Ӧ������Y�ΐ2��q(nbkj�E'��u�۬8Ҭ�vk���Z���eCH�12g|ٳ=�[�d���5��枯.疲 ��Y٧��
�U#�;Sr���\��`�>[�9+4�tr��&��׃z.hgR�t]S%ZH���y����m���{@ǖ�Ymp�����C���g{r� ��-vצ�4���p�,YJ��WVV�g>)��yTPv[�G ���E!? }+n�	��CL�h�T��	�="@ࣾ��d�_�jr�׺c-XN$<1��,���oe�jN��VY}�Bm�>m�񌍄������[�n���#~� ��8iMWW����B@Ҡ�μ���W����C� X������+m��ʱ%�$��j?Ȝ�ǳ�,2;kM#|�kW#w?��<��V�Y;?>�$K��K&$_R�\b�a��@$~���h+t�,�R#��I��L�?[�pa��ּ�@t)��u]]��7��I	�|�w�|�A��ۉ I �	H�E �A�ˮz�h������ߏ�	����O�/�?$NX[��V��"9�͗���H�kEz~o( Q�+o��v��?����,c^��?�Ǌy�� UV1�e�8�#1J�1�C�"���s̻�:׽���U���6s4p���/{V6�#����^nK����L��zר���tf�iM��H��9��/4�H1r�C.���,�qH���A���Q�n�{լ^m}�xsL΅��������~��'�AMM�����ߛ6"FuA�άG���	 ����eke�	��&�-w�n'�.��8Ng֠&#P0ۊ�����9 �^����E�KA�h�:����Z�wh���u�JA�zΧ���+���R,�AY����j������^�*<���y,L�z���(}�Ǐދ���K��O�`y��I/���]r&6�y�	��a2�W�;��+ ���HMRH�ߝ��#@D|gz��f�QIN>&����ׯv���}}}�hYAn�Z�۫;3�H
Sָ�*L:��ZU"�e���hr�^�t�����Z[[�tae���>j�t������r��5!�޼c��o�5=27��=��z�σGF �T��(���� �d�&��&A9�	�e�<��D$�.*hC@���iX��J�m�z�v4r����j~7FJ�3<���ێ???t�X]��K�j[��n��W�����q�I��>���@Y#[q�:�B��_;{Wv�t�G�h��Pu`ѠZ$�31!�#�}��٢�39��V�"Vؚ�����:��DL��_�D�;˖;�[�Kʰ�KC����\W������<��с��y�grJ�|��b!;[���h��	�k��F�Y�*������ڣ��5%C����������>z�SU��ڠ�������\jQ̈��:����Lz��(�wJ��|M�j� �Č�TTۅyP�a)�b�ͮ
�t�:���<�j�I'W ���L�vy1��Lҥrsmqd�t���!����k���I�\�JF�+�n}1��k]�������9 ��q5��������n�K�X����i�<�������V���k�G(�a(]������ˌl�T>�cC�-����q�lq_r�,˨~8
OP�V�Dz�����q���l-���n��֕�f��\|^:��<������D�:���w�o.Q�}���4��d@ܬ������V����f.3f�>�N����59R�E;�e#��={��G^�����-�k��˃^���Hw�W�������JO/$xÒƹ<+uU��	pjk�/ScE�b����
Tf%b�s�I�8��0]�P�zXU`������}wJr�򨚯�Qn�XY��C��� b77�d�z�5���jY4�0��v�`���T�?3�.�>�[���(��;���!#���k��������&F�#n�<p��Z1��Dt��I�[���Ĩ������n���٠Sc�cH���r�� �^��+�e
�]r�H\�ޤ�P@�ʓ�z@NU {�#ĉcχ�Ţ�%�I<��F�5�d��unG{��>�� �����?��h&��Uy�iG�;��A��Z�j��S�u=>�[R�Tz�AK�54�lW�J?�0-�DNN.T@w��Y�WHHH+��sP����g$�t�(�����Aծ�E�֛��*6�sC#�>����4ͤ��b2��U��RFq�!f��qa$�Z��tУ�p$�M$yPo���>}���d�e�"� �����
����~���5�������wY��lm������P��;�H3��֦�E���2���#�~]�i!B/ڷ��5� ���>���붵^Z�7!v}�{2��\���x�@"�!:%L��ub����u�u����uS�_�
w�[�UC/&,���M�F�[qj�[��X�J���xk
����BY���LAh�;(m:�e�uV�K�L/Z��ͷ�<-����[_U`?5�F�U	�W)�� p,�����O勊��'��Ļ�t��;Q7y'�ꌤڙ�9����;�Nv}1��Z�(+~�%%rF���^;p���bSp��a>^�������E�|�"'�豍�a�H!B�N�.��T�9*z�<�p����^�J%��;	nq��	A~Ѕ���A�2 �k��?,~�i�y�瓈����4�/\ �v��#GR��LEDDN�5km�@�P��Q�^�=�D-�i���3LXA�9�/��摪)�Zjš�r����9= ��G�|�y��2��y� �����S��?�u�`Xp6`�C�M�yT���\Y/5����J�e������T���Er5���	�_'m}�@�=#�Y=����j{���݄LMM��(vD����A�w�fK6�Z�-6��S���l�{]n�8��2 �d�����[�0Z���5!5X/-�1���=lK���xB���h}(��Nr��w�a��L4@Q,q�a����6�АK@#�~�n�\��C��;,�;Q��~���Ym�O���d�����ٖ$5�wg?|�pu ��DN��H���5,��U����,�VE�Z����h�'�ק��w�%��)Q����FM��d��ڸ�:t(��
bQ
h)�)������h��tu���wf��Pe�&B���윜�jRo�7�*�p��E�|UJ�Tv���J����e�xOy���	4��}���d�1Dj�ȗ[ A���@1
 ��H*+5����g�Og*5�^��X+9��ZT�@�6�)�z'em,::w�xV�I�7�E>��.�?���yk��.j��]�0��SO뽈x�����)Ӽ+�(�RQ��F>z�������*�4�� �! ��L.���e�mq�1�&E�I,��&5Ŀ�b9~���*�D�qMwe�7��]1��ƥ6��(5�\���%��H�$#��/�U�Eͮ7�[�E��j��o��� h��������QSG�}� sw�h���i+~i 㩊�E�<�_�Q�C�7K��R�&��{
L"�C�\_ڔi|B�l��;n�<Y]����)����=�)�������� o�l��л�4�=()ޯ[ln��ڢ�GA:��>8ை]sV�V��QC����?���Ċ��A�M�aq�*���D�����6�p�^{,ڽD�|#A`�V���h0��!��� /���R�C�I_�<$X�{EEw���5g���t��󽣣��p��WQ����މ��$>���M��8a�k��dv���t��>~3�6(ҫظ��������V���-���^ۦ�9۫^��h�BK���.���R"Ov��	�UV�V�M� ��x���PTh��.��L���0*�pr�zk�T���Ս�mw�~�EAH0���H�*�Z��3$�;!C�W�-)�$��^E�L��X������ר�[/��kb����4��9(YyUm��O�B��I8Vp���]��j����aU<AD�α=�`V�b����Ћ�f�p��,@�RL^s�E5�. &�J�kf���b ���ב�D�vB*Ǡ�ɷ��蕀'�gO8��a����r��'��2n<_6��-4q��@	�Ocd��X��dJ��E���|m`_l9 On�k�72����o��3/���|x聐�f�$�-���@q�0�.���Ҙ$_��ۍ��P?�� -�EcR��_����lm3�*CuS��zvEu�N� �I� �Cc!oI��"�1=�W��w\�&l�g��P�+E(��g������Оj+�; �"׊�� ���=N�\�m!0�	���bI�1T?S�Q� �i_b:_	�R����!�$�J�X�e���e��9h��ѣ�]��);�~�8\#�mM<*q�7�=N�oh��_Z�L��l�K�E ��W�F��k${�����Vl2]�e:�@�_F��J�����x3�N�3��ه-�<��ޭy[�a��sL�XE���:ț��r�GιooBE�z������qa@;tF������B����������x�D'��I�>�o�mm	Q�f��A�9+4/��m;�y�f���4�G��j����)�趵);�Il�+I�=���>��=n�<&O�N����E�j�1_6{*V�갵I�]�����rJ6�񗶳�Y��,u����vo	%����R���N�֭r-�t��_ZZ
�O���ܿ��[�6ٖ��חƩ�=�L˼��`려�\h��襊��#�?��ff;zzR�����Z'''-��h�>��H���n:�C�*�ܖ��Os���P���~�����&��/�s@��\K?���#셳�q��bX����vM'Ǽ��!&ZJ�ߧM&�n'�F�c!�2}X�e�;!J�-��Fpj��u�:2�Ęϳ<҃�����/ `
�p����&��Fb� ۾��Q |N�������;K���w������G��U��+ߗ�LG�ǃ�n�|5᭳��Jͻ�֍�8���٩�L�ۅ��&x�^���饹RQQq�ر�,�7o�����v9��݃��ۡ�]��/����Qx��~�o$a��cC3�*ڝ�@o��a)p�"D�k����bI!z�*��b��ddy�uMS�u���e%��&OP�N��7a�O����h�q����vQuuu�
�5E�"�͟�mKz::�k�����)��G��Gx����yH�:���n~�"�vpZr��P6�Q�%U���$K\����ӊ硽�����j��;��;���qff�<�6b�ODJ�vۑs�ޫ��u&Q���s�%�4ѝ�@��#8o��f'�ޗ�'ޗoQ
��(�����",�1��-�~�����?5SO�t��c����X�ԫ��jI-��A��%�E����\�����GI	�B�S�Rx�B����5�����#I��N�|Sk��=������Xj���O#U*�*���2��b\�V��#k�y��1�1 �A��_,�$�P?\�JP��]891�^:���������X+��}}6K�RS�鍞�"�YZB�ûwe�yo�T��b5�8��76�)R��O�{Q�h��yT��E���?�NX�^�܋�Ⱦ����o�1A\]]9�Ѵ�8P����(ٻw/tRc��w��sk�o�魭��R�R�� �gclgw�T����sw �d�y�����޽V���^�u���Rn��ȑ�A<z��� �	}�m}�f��(>�3o��;����&v�Jw��������T�q����h.H5��fѼHYQ牗c�� C�l�-��^X���}��L,B��ho.�;����uv&�1]0��=��y���^��[����qϞ|��R����}�����ۄ�)ja*
�']yF�떏��׵>��>�m5l�wԤ�_��~ǂ�4�f8�]~�Ǐ�q��iR�9n�,�>/..��eb��c�e#?U�:�Q�p.T�Y�[-�tttK)[�Ț��"��=g7Ǩ��W�SsC�
q��6~~�켽66&~Zex�ɴ,{�a�$c�&`ju~Ļf�VbIZL,Y����IST�� Өك��^��+w�F>��?��q�>lq�i*�t�SpX����Nɬ�b�zK6ߐ����������{�
��%�SRlul�Y)��Ś�W�,�d�CN�� �M�Q���M�U�6����<���~�G��I����d�j�xzRi��$!�*+_LP�l���u���I�����U1^�=��bK��_����n�w
����m������zP*$���S5�*������sL���JC��/Z��=~��6�?[+M���;�[�5�VD���s�,��\B�/g�<#�^b;���}M1��p�����0��	r�llIV�'�M\�?f��t5�ʷ�vnw
:�"ǑV��������$C��ѓ�2鋏H��-=Ye�l���n�u��Լ�˼����V���$J6iK	�:�&� aR��e���3�;������G�F棄Ŧ�,��#*yd����+�NQ�0e�iG}����9�B_��|��K�鹊�v�ޣ�A���t�\}߅���Hvm�Iܖԋ1Vmg�ϱ�v�wgq�諱���&T��S6�������q (Z����(��;�Q��Sh��1���F���-4���_YC9�����@����S��^^e��� b4�{��ڰ{}aBJ�ݮ��H�+�t���F��2H����I]<p��wX/�̶�$��mg����s��u�Pb��SG��Р=�kn��Jqk4"���NC��/mO�yԥ�{��2��,eU׻� ��g�=u��o^i'���(dD��y�@� .��_�|�p�&���ƞ�}-3DpC&�-Z���$}}K0�����U�`����FNP`b�.�#���?�rnwT ��;�G���4Y�E�Zo��"��܏��|�:ݕ4>O�x�VHU��l� iY�997?�ja�� ��6�A�C�[���=m�2�g�������R����̭�k�Y˼�=������˨E��̀�5�\�T�Gno���j�y���/v����\Dc�����K{���cgƆ�?�����/P��R��x�}�)��2t��auhs��b��^Z�!Cf�tw�v�_C��H�2��>1���;�!*t�aO��۷���i��u�|��bGc*�_�����I~�����__'�=-Aa�Q}鍴�FU��{�T�)�e��&۠���)~�JP6�q���5��5���'�R;�̐"!�WN���>9y�7ʘۢ����T����I8{Q���Þ��t��3�ʡ�,d�o���R���(�����t�����^#�>h�qw�_;K��?�-�6��҄oR:�]R �5@b�����y�"����+���4jz�1(1�1q�== \&{�5��<#��i�r���zO豚��g��U�|���V�%#�mjgx�}��)�!��Z��8Q)N����c^���x�`��tCȘ�:�3��
 9�v��{�'��j����s��A��S�Ô����2���2򙠐��)r�$�$����>S������DL%��K_��E������K��z�i�O!cD^�����K��d[�(�_���C�[���Ƽ9<�w3C��&V#[J(Đ���ݒ��W��.m�d������J�tcy]0�HU�_9�zH^��ڏ���C}
��"&�n~���;�6	�P���Rw��+�_e��۫�ٞ��������q.�l!�0t���p�~��*ض?#Gue��2��������Ae�E�p���cC�w[G���H{��+��
�w�1�A[w��ȅfk�����HGIE�nLMMϱı��_���&\?����b��a��]���Q�o�
��1w��a;��+]x翋\O��UK�>�\סֆy���g̏���B$��{�d�~����+�d{����cQ�t�pxOz3�3=��r��Y|�!�m�T��oY�t.�������������l���A��W���fO:����(���r��S��w��*)K4�AK� �������8,b�y9&��9�T^߬u�.�;�M��	�j��F�z���$��^�q�1_vO
g!�)"`A|85���65-�/0�)�]mz�Չ��i:��|7?����BY���m����+-�}���!!!AJ�ݳ���"0�/�E�Ӊe�a`�^\G����{r	����sM�@,#<�0k��� ���Ni���Q��A^�Cd8�x[�����mJ��eB��ݲE�g�R�/=�����0y���s�K'����蔸�+6��ʹ�B�ύc�ȋ�E�9W�Cd�&�%	ꮮŤ�U��:�Wh�_ؕ�8bq�������ْ�c���m�]�R���+����!:����XyRB�u�q��Wm��������^jg��S���v���[!	jn�Yg��h廒�M;s���:>a�|��������vtdq��t�x�v+�����7b;I���JoM�-3|mu����&9�!r�n�����o� #�LX�Zɏ�����-�.�BtZ��kQ���G��n�-}#��A��!J�Mnz����X!C�&��]��{N�&����b<��;19�˟ER�&���6�x��)��!�hB8z����rG�¯c,���, �4h>h���iM.�I[�����^H��oG�J���K�Xp/�j�V�,�BL���*\K�.O/sh�ݵ��u#v�ى�\}�hHc@��b|.�P�+E�)0|����1p8��꽜�詺o�q(2�x(����uO��?���^}-����Z*�9��c���7��fgg�t��鯚��Q������j��ח>�����Y`��x���}�(����]��~\ϟ���ŘE�r��_��.�.���{g���K�QFSS}lC�߀A3:����>�N�w�7φ����=-�3q�<Gj�~����Ò̀��:���O7���K�!i�U��Z�ka�����ho�٢�.
�ٸ����;��w�k���
�k�����>�,�'�6��<��[������'��
qο�(�zɩ(�J��YS��XOAt�7I���%���*�J-#�݅�<ä���%ksRL�:̶����.s����������ʇ���\�}���/�R�]�)\�z�N'�"��gOP:�8�5�]���<�|EED��/Q�w*J/���,��(�<hf�.|�8趋aN�_�(�/�ɲ���� �|��LOn�"�[�V;[+f-���16�Sf�ǟ�y�S�Z5��$�tT����<���	'�[��S#m�աW�6�W[4��AҥY�*�$�b�ݐ�ӓ���2�Cp�*:��Z��W��!j�w�X~�Z+� f��B�b�d]�jx2"��Z�)=] >z袏j0�/��_�����㠽誽MJ�w'��4T��7@��򬒯My$C�%"��5\���a�4ٖ�ݕ�&�2t �t�����ҭ�RME�W<�o�ȹ/^p��L����1�8C�%����g��u��S*��³��%[3�f�o9atʪk�������fpG]���8�@��ig��y"!T��b0ū��I�ҏ�f��wc���IM~{��kO�B����}���.���:���nJl��Z����]���[6oUկE��y6↬�:���[�懫 ���i|�,{��5��$�S4!�l5�x�ڒeT�=��mS�'n��!��B�J])�s���l���M���o�����e�?����\ �J�_��,2M�*�[�ы�餜9�8���+����I�o��Q;�@HD��z~1J]ye�*��9:�ݘ��[gѫ�%qz�v�7��$ ��t"Nb��t<=�t{��&�l��=�pʜ�r�Y�~�����ˌF�ڣ��t�QEy�2���tT���Ο��<�{�C�EE��h�V]樜����ڬ2���W�k�]�s+�=���uE����k�6\��:C���>ɝL�gձ�ٷ�	/���_?K��hk���(��m���[S32.����"���}��制�����̫	o'�$�`aa�ε����D���{K��x�{_�`?�Wޖ|��Qx�T���.���Soj)�l�8�O�+����cm����1'�;�\���\�&��:��b���8ϕ���1zkڄ��&�6�m�*��C��g�������V^ZZB_�KE�T��ZZ�k0�Rc���#^^6|�i�r���8��ӧr	Ïy�)�xw4�3��Ѣ�=~)?e-�$ߣ{��Y�Lu).����4K����%+�NJ�e�6���2j��K��J1����3�L���%(_�=s����6av[u`�ѡu`�R�j�t��E3P%���C����Fi/��+�R�������i������.TL��i��<o��yxk�׏:Ց�o�HС��˙�n��Uǻ�u�0��]�堂�'���GNĘ��#��cQ�Î�����"�v���4aWƗ{,/��u�50�4�ѿb77x�E��Y@��ޱ��S�}K�X8���@D<厫��G.�����(����%e�W��4���f����D�5�z�ޟk*A���͕qe����n�1��@���ev�L�|Ew��>T� iS��[ink������))Jm[��-$(1�Bf�82��:�뫿�IkP�ů��W�{���'��`\�%��
"���%DE\2�R�|������s��cLZ�n���-H�|�Qp�	z���.�|��e���W��]`�X�rrB���j����C�#u�rY��OR��R�?w���<�_�э�~u)��l����F�_����v�>���,\a�)�9�)�}Y��s������c���S���B	�O��ו�Q�E�F�g�KC���S 4d6+d�7vJ�G0�!䏱�ٵ\�zWM�~����6Y�]!�_��[)��b��x/ھa����?����c�KE���[���W���%W�gd�]@��C'�Q�QR%��T�з$I/���̬�����
�h@M<X�r޿5�P��yK�e�QLZ�5j���H� 
h�ɥ�`cj}��Au�+��d�P��[���j�4����l_Q�?�2��e1t>�[�1~Y�o�$�T�:QBQ�M�L|�׶i�%�~��QTt���+%+�HI�F�S��C,�����{����E����-�C��!]��^�Yaz�k_������zS��n!i�>��t����	WEw�d����	$i�2�qV��,�_t�/0,6J����z�_9W�?�GK�P���C憸=������N��^��d�J�dd�D|
��q;�Ba�.��%}����-��9o����@���WJw�-Mch��&2�@�Z4�D�.ko�9�7y���c�)=�f�WL�ج7��GE���9[U��ۏdTx��B3��'��\�awx6%>��a��k���z�p۝���x�iJ1�yX��� *�ƱmyJf��������X�,�V2���{��*C j�YԊ�c�Z��\�۩]Ob�\����[�O�|�2÷�2�,Ym=��$Lc<�kL�M���W0VU�Ϡa�w�ng�v"��	����Ɉ�k��.�$��.�=Du̸'Ǣd�ɜ��ٝt����"2퓀�{�}�#~*G0<:Ntv�����O�����D$�d%[���{��I6%�Y�:6ǖ�G��=��:F��{?���z�����k�������q�E�]T�q���\�w�,"Y{�)W��u�f��M57��߳5��7͛-	F���A�0��D�L�)��6ً���V>��.�4PX.t�P�5�J��P��-2��Vɿ�@?YƆ�n�m���Kj��ܐ����ż�\��G7M�nr�s%uNņ��-ٳ��3�	?!�͋!1ʿ
��u��Q�_�ǵfj�ʹ����izЗ���%���
��b$�p�\ZRR��v����9�I2�
r��ouU��-�r�II��|Omȧ�4��_��0���t ����p�}�!�`�����*|���:�ai����߉����0<Խ]�GǺ�U�Yҍ�� �����C��&��1�(���j%�B*��6���[{'3��;�F+.��0}5ͽ�-��1���dw�=�IC�$�c�50>>؆���3�gg��ɠ��z�ʦ4�u�||�I���ȧ�<�U:���+�X�o0,��I����p��학ÚM�PRX��Mӯ��օ�;~�􄉍�do��0?ez��3*w�2^���a�
	�e[���j)�ll�G׶f����-@��#���Da)�HW9N�s��~��P�M�{�C+;�V�a�#u�G�6�*l:���Dǣ��m���pd+�w�u���?=�>�k�U Sv����^n*���t�ı1��t/L����Ģ".xgV ���c7B�[�U��@�v4��F�>i������TC
���gL�~�ˋ�÷���,.�KXg�z��~U�%/�1��9�c�BČ�5��(��M����U��}�M�%,")S���+���L���lS<����	:6��|��`
�F-"ј�B@@ *����=����������e�%��/�����]�UWWw0Mu���q���NIĉ1PU�t,|�6��G��zP����~���v��z����r)�X��*e���E�]*�3�>,�UB,-E��%�����o��{��fCC��ȕ��·+j���P�q�Y/�j�����Y���8�p�q��E�m%����$Ac�x��t�q__��8���
��SgE�oH�/iJP�/��eq�&�=]�4���~4s�V ��g/ˀ��$����	�e;/��Y���@����8�jA�"��zF���M�����U�a:�M����G�Y�A,�^˚a��8j�[�O�%ʾ��tA&�~ˍ�PQ��:�#��ԲL�o���`��@��c����͌9��ڽ?>\Rd�hd��ʂ�+�,F���j��g��c���(��<-�mE�E��
P"2@�s�%���F����78���us�9�k�:��߳~�$�'c�T�hѥ&�{�i��q@��A�*�d� 4р���;��3r��k�j��=�}p���=�-�IFVV���`�s���v�A�J/���gÐ[]�n��_�W+4	�2�Cb�s5�D�}�@�I�eڷY�<��{19G?p�OntO�r��a�tl�m-�Vn43���]7�x��I[$'�(���TR�9��j�j��{X�	�VI���Q(���r/���6C�� +%������ɺO�ջN��Y����-���Z������EkdgZ(?Iq)��n$eͣ|3�oۜ�Ya��[͎�9/�7��Y)	���E��-a��""ȣ=kx�OW�����'��0��R�'t�²�Ӵ�U$by��"���ox{�Ҙ�Ş��l^AZ�y��T������R�ɩ<��j��A���4��F���z���+ϔ��OP�2狤��K�l��y�>Jo����d� ��i
&�
� �K��Z�b�:��Gӷ��1V���F$��>�������![�]�)��b�c̓��K/�/�l����L���>|8�(`����BB�)(�O89�
�]nĻ@'�3��c���<����D>6Kc������>v4�cn*��:�v������J�*�$�Js�Uv;˪`+�!���6,��і�x�^�.�LM34��jf�@,���o޼�"�/ ���Y����G��0?0��{�!M�gʲ�>Ii�N��3��@π&&&)S�{Ƿ�&�J��w1B�<��%��.ح������޷R8����T=j��������||��x��5���0�ۼ��S��fJ�2��;{��rU$��[���ȅ����r]o��N�k4�>2��k��`\*���	I��L�7�Wy�͞e�9��~��AZ�(
a��V���3�0j��O��XH��G�Oa!R��y�Ϲ���J�a�w��]L���՝����P�mʞ&�aǗZJ��3X����(�[���1����] �g82ן��:��	�ۖ�wT'�����>ۇ�>ɭ����G4qU��?N����^�^�M�s[�}B���*���]�$ ~A�w������Ӿ��B�H�HNdČrZ�4���1�
��BP����''nJ��[�o��,JA}MyL/�h8+D�K֜'<�;fA�*�#쿇���(�ei��C��p����1�aW)��?#�%E.@�Y�H��c{&v2k醰&�_(��9�������t?ΓhW������%k�D=|��G� ���2������̃jl��Չ��w�@A��3�U�rF;�>zx��7����Yk|���wZ���t�\w
����$)���m�+��&PB,�>�͏B�\6=��=O�>���p	��%���%��O�LC��ޙ���;�o��<�OّZ���m�?[���JS �WJ�}@\��t�׊��3�´���N��iƁ2�~8;���[}B��}�eJ���睙��!=��4��%r8��A���U)�l�W�9���W ����'�DQ��=i�{�����K�ǂdr��]������������7��m^�>�M7:L�8�� �[��䄠|��\{W�L�ś�*Y4r@������D���v�~�����c���`���$b�x�Fi>"4!A�#����->k���Oo��@���� ���}_����$��.rC��Z�=3h���ʇW�9ov�A�g�Щ2��|gG?��\���}�>�O�������"U���&�W���+bMA���OC"OJi�qHe&k��I�����-����*'V�9�����
4���bA%�������~����m�Q����zyݏ$r/&�����+�.}��<�����{��ԄS%�Xy�[���Z<�)nѲJ8$�"�$�5��H�� ���կ���w�at��D.��1[\>o#�귉)�͇�Y_��hX�dv��¯�ZO\�~�r�)���׹l�i�EzM�ЁAsg�e��v� �P��<�<&�@��<�����Yo���[��y�2��G�]���'�$丽�˴'�a���52`�wC�SЛ���Ŀ�)����7�,+�K��l���;ޓ$��NXsUR��B{G�B�8þ�py�Q�XՓ����+1|�k��L������L�y�*�����?�-�x�'�sQ-���{r�7fM[c;�3;��$6���(d����[r[=IV�����n�^M�?��%W���������ܩ���!eI
�i¢��%z��o-їթ���?�d~0�O�>&Ƽq�~)�N=}oC� �#��fK���r&�{�I_g^�㩮�N��TҘ��j'-�S'F��p�#�d�y�m@_��C�hsgM?��_��_Nm����7k�tZzbi�*$z.)8MR'�1�}��c7dw��G�Q��I�@R�����pֆ�7�s�ؠ�R��S��ڝ�W��S*�z�2�����"��#����+jr�������%�Zʗ�Q
==օ3�0�=�=�s����Ŷ�J�Q���m;�{:kJ����6��f+**��V��p���g��D��X�v��fժ�%��u��ϔJ��=��!ї!o��{�p���z�=IcM�<@���f���deփi�;˚�R�C�|�t�H0�ޔW�K����-[��wlo�h�M�3��l%>N����u�N��4��k8e�M��=��}��>4j �35A���?:�Ps���`��[2f�h�+yLE��@%�iC��+{z�񪘕����Ċ�M�ɳ��yZR��n1���yz��}u�^�k~���o�W��s�
�ڲ�Y9�N������vS��'�=�I�&��3rvR7�	���a�BP�����Z�($�����!���U��$r��>�فW4�!���RN��j9�iB8Ƹ�[�(�������k�}&�猷]P��]}�?�j?����+N���@z�?Ro�8���h�GW�^H6C3+�D6q)D)�8l�A�Ɣ>C�m��i�-�1�
jQ�x�r٪�ވNw�$�%�q!-��˟�G�ǹ���L�d^�Ir����d�OԤ_9M�}
7�ξ͙�����>GN����􉲖 �W��D��E��2?�K�!e?�^!�Ξ}�T��|���jD�~��a*\�J�n@o�
��Q��x��J��*�@������S�L�5!anV��S�ɉs%���򞑦��Hx�"5���m�W�u�� �<�`�v2�D-��c��?b�
����f���b��_I��+�~����V�zTڎ�5Y?�ʩ�T��$����Lٞu��lE􌤋�0�.��@�W4+�άYQL��o�%^w�z�OÕv����T�`c�m/��p�.���OI��'�- S��	"���i�Ib�:��pP��KN���LH5@�-�����bE��͌D��B�m�x.����~��_K2��G�vS����E�๱^�M�<�19d�TaC<�E����,c�g���4�Y<���h\����m�v4x̾�?��R8�P6ܵ�L�?��oXCٿ8J��l��#�:��ure������fM�[4~8�u�L���OӸU��O+V�9�J�i�{�z�%w��㉴��ZO:s$�X��˿�0fc5-J"@.�ݬ�R�K���;�Ig\ϼ��ÖO?=�{�a��AP��KwGUcN�ꃸ.���֌�63tz/��R���'����,M��PD�(�*w���
1x��yM�]Rƽ�x1�S:~g`����������T�l��mƼ"��Fwf��}_���CG�}jMi̝�*��ڝ�O�Y-5�O��E����T�2�\e��D+�e�p*�m��H�7ۨ�n�i�g��)��;�$�ʘN��h[}Y�ߨ��HRX�rzٶ��6�ۡB������[��ؑ����I�7����5��[��@ۻ����o��ce��gH�p:MKrĘQN���몧�Bz����]jN����$��q�S�Y�����7M���cNZ����cUڤ�b \ ��6�n$�Q�I�0��b5��R1U��� �!��`�LO����νC�4Y?��\dTC~��/lf~��5B��*?V�L�i�wQ��1^ާ��t�N��[�;�{�mkH�h*��<�?�!Y^�,�#nP�u�O%}��>C�������K�zi�+�i��!�:��:�a�)�2:���
�؟K'���)���I����gWPJLv�}s��qL�T�>�$���!��eX���n�+V���H�*Nek9̥*��׺��Y!��t?���i@]����D�W|v
N��k�$[�Ѩ��[��רu[���zE��1B�<��W�:�{ʴb�@�9a#1�D+�k�"�h��"��?�>z�;1���4Lvj2L ѿ5b�Տ7�Wݏo�A��(܍A���Ӏ����ϸ�ֺ��%G�W7#�'������Ahb��M�\Ţ!v��Ia��ORٓ�����9'lKL��m��#�c�<ǲ��1EA��o=)/-2�P9�D�D��/�x�	oN���x9L�/eZ����,�sJ�I��i=�����y�CWr�O�-P�rO��d�F��s�Dt�/4�\��������ԣ����[(��E�4m#������p���b%��Jsv)�x!Zq�"?r�+-�R�����\wjǜT:��7�SN�#��L�����k�@�Z8u2s�+�@=خ*E{�m�����O"��� ��ܯ�k ����.)#p�
B�ib�^�T�#2a0�6�a�=Q��d����+�R7skM������]��/�-��x�秤C���y^���E��e�[T{�L��<s.%���n	��k�?N�?t���!RD�^#9�N����*���%^����'��\eZ��e����������}�I#��#�)}�qJF7K�MrI�b��Ӓ��3Dgty�?A6��|��aҲl	Q'��3r�|�^�x3��[�����ؽ;T}Ya�lT�Q�2�i��*�����W8�U>��9�w&�L�跛��7z��E�
��G�MI�Y #�s[+d�43��\�By�o���LTCG�guB2=#B���o	r�骸O�2�
\�I&"B�𱳴������@�!�������6 4���5�;_�{�KW���_}c���ڧ����P*E"��x-��H�򶛼��E�W���{z�C������kr"�ْ�N-�g�����=�4��)���o�@lC�2=A�P�%���~��e{L��_��ڗ�;�U
�	��D��.�'f�,�k\T�	&�����H.��N�=m����������X��T����'�z�kr2[5��LsyrkU�es���.B2o���f���m��Q��8)��վTJ�����0ܿ-��!��ju+U���E�%D.J6tTq��Z�S/�D],��۞z�e|���ﭦ;JV)u�a ���:CR��((�G9��z��o��摪}�Bi�i����A�.DGu.�dfa1cߘt����c�����~����+��]�
����Y���7	1:���!��1B+�!��se�'�631��d��7Y�Zg.�?�=].k᫉��� ��Na���\ʘ���oٿ��9D<zQ�`�P=V�-쇳3~	����d��S��˟$�p� �8_S�9ɣv����k��Y��h��L �C��:��w��0��v,l��Vjq#�U~�e��<�$-cɜUk7��7|i'o7o ��fg]1/�%koS���H�����Z*g�����-�[�� iG&��!w���mD@Kea��.V�C�Ws�+�{��������g���?Dh=MV����L�J;��a�g 5��N�ћM5�"�
M�Fs��A��N�S�yw�]��@��B 5���^�?��\�m��jP�ӷ�N7m/NT�4�;CPn���᭗\�?���[;,s5؉ۅ�ǖ)??�;�]����ή�c��t������J7^�$�%��So/q*��u�ޮ�~i�,��{�T;��~�-����%��7�h����w�L_�_�U� u;��FE��X�mۙ��-{�*���J#����rB|���=^�TLcold�|5��n5怏2�mI�8s5�D^��i
�qUC���dW֬�O�[���K��g9�E���<�>�'a���l�F����ơ�Gهz�2�F�mf{B��t2��r��eS�uW��q�٥��Үu���B��詡--��"],�HB�و9@�5�M��c�z��"G���۲��-�u��\ʫ�vvb�6�|�F��.�B�H����nx�z�ZQ`p=ܢU�E"���|*��-������M2����.s8�$le����1��P�Z��+�>(^���¶|sI�r1��c�5���ǜ:c�e[��/m�ɮ�TEQܧе�Qz���_���:S��~1o�)���&��_-���f'�)m�.�ӞFZ�}����S}u���eِϾ���إ6��0z���8��x�C=3�v�l���7��M�f��A�7Q��;
��|"��d����uj�5i���__Y��D]rD�|�s��W���Q��ߔ�6������(Ʋ�:
�� �y��?�*�YP���D1�&N��H���/��;�i�=9n	k��F:�o�,uv=��{��Y�k����q�kt=�Uܕɞ���~��.b'�5Ux�Q��ѭb���Y�t��Kɰ`ݻz������1���?�[L12+I�QQ������D�?I*]�-��"K�����az	z�s�q�u��.-R���H��a������1��1`���_�����n&io��>3>Ԥ̼3 �/$@�u:�z��5lr��ɥ�'U����6&��Jh��L��e�/%-!����4!�E�q�ƴh�	u����K?FP�<���ɮQ���mc<��[x�=�;�FT�ɒ,_���i����(�����W4\��R�7�k�?�b}�}��Q�c�uѸ���!��ܧ�3q�I⠽��}��u�9�E��G��!N�ؤً��>7}I�����d;�޻O(�X��:�9V{SMi�-Mo�Rf�v���t
ً�����΢f��8�I)�#
�%�ªv��0,Rg� Dx���u[�E[���YH<�|�Ƙ>��ч�a#���c��ƒ(J�/eÝ�����*��`��1��ot
���宋U������'^�b 'S���N�(&�UF	r�1Ug�\^R��|)af_���+Δ�1ݼ+�����׋��d����� ��}Ji��X�����O*���P]R��X�7�`�g���xՋt��������fk�T�0
�CO��#/���݇+|�}UG�P��G;�M�D=W��(�W�46�$��o����gP���*&�1���T�Y5rD��!�*��i|a®���-��񮾔�?�}_u{zTO�
�� _�ք�v�%H�[�0��Κ3�� wUrLE,���e~�$�
�-��^<���RJƥu�/
�}�mrү6����:]��k�Q�q�T!��?��TNK�Y���3]��E��H�=H�W�})��4���?��F�*�
D)ڪ��!p%��U�Ēv��mL��=͕�;]ߖ2���'�m�5,Us���V�I��Ad\�+���[?�>�h�n~��/�m�e驩D��j�R�,[�%�砚���ᩎ�!�t�T��ea�C���wr�XZ���������U�p35<h�&>2�kH��W����;�����>������&��8V(�����Q�����E�t;+o�n�<�P���Sea��Q���b;�Y ��˜��u�s�y�sD��`��}�fP��2"�+�3��]C��LTC;>b��vN�^5:���0.Le�Ax�q|az�N�v���1e �⟱o���,YԿ�\�,x���u� Mpo���_�4�U,�f�X9�5[�>|�{��nT�u���Vb�NLذtfJ=Е}Ԉ��+��]m�1YA���|�}��a�ӑ<��,�{��dl|�}_敂]<s+�=2��/!ު����v��*�����(��EU���1��MQ�1�nYL�ë��wr��<J��ƣ��[���(��1���',>�9��7�o��q�U16v����m�@��Um�+�>ʅ;Ց/������&٥��9.R�~��Qĸ�E�vl�)��G�3�`���߲]�e��MeyWY�v�֌�g��kԧ�T΍��T�+G�����9�+G�A�2H́�	2��]�n��ۡ�Ud�����
�����p];�j������yD�uW<��R~(�l�d)C%]��(t��-�~8���c���U�
��pVZ��雅!;���ƫ�/x�Z��t,B{x��N&�v,Wpi@�	�8���[Jж��!��m'%�۵���6�>�!��R���&Bn��uƻ�Mc�i�_�W����Ϣ��o4 !t��iEZ��i�|g�zy�R��e3����[�i��k�� 3$x�TpXv�?4o�h_��:J�8�NYu=V��'
;����ĸ��ҿ�YWo������R�O�[�>E�e�EY�a~6�Y9�5����o�e�8������y�	C�\�8�x�ѡ����ÍY��CJ9���� �x��!�L���mm��|�<���sW\ܙ	ǍE��h�|3��C��F!h����xu�ЋW���k69�:۞��Ē-){J��8�@w۹'�"˄��z�ʧAm����F_���ŉ6��j�-MvuAz���Od?5��|I�ѣ��:��
�y����?� �"�fۉ�P�ӭ�^9S���ue���Ly��n<�K��&��Ŗ�f/����S��G�AP��B[��Ѯ%)��A���MW����H�{���@?_���q��]<C�Iٍ�N9����RX>�9���e;"֏��J��}� ۏ�jLe�t���	�V�l�(.�e���x���#ˤ:8��/}XS�Ȟ^���hv��mҺXͥ%�^ 6!k�/��.U�+c�D��]�\�5��UCC�E�s
��%G�6FCn�z����!	�����9gcv��mM�5���羉R���]��u�r?'�{>6މQ�K3����8:�c���MR���(��!�5�Z��T�縛A�e��{���޳	D涓�lf��&c�
��҈W�u��H�؟��/���k�yzAy�N�F�(�%�h�q���Ѐ���C�CM�;j>�9�<.��OO�pwa�����e�f&;}����͎���\^5����, d�
J�
��JΝ��͵�{s�)�����|H��? ��طy�����Y����$3V�0t~2?�q��j)|=��&��\��O�_;�BqWo��gF{��؀�*1M_��c{GSN�:	���`��&������07�����n1K[���m�i��k�v���F������dO�l��ӎ`���N��P��.@�R��`�$q��{d�b�1��q���Bl���~�SEcK	sP��L1_��"� H�N�rj����<9^v���ތ8?�����o��h�r�8��
�.�Κ�V곊���?�vǼC'F�o��䎌u��O�:�6V�U�m�I��0�|S	#75��,�+�/�H�y�6,�Ūa� :5�Oo-uz�������&�,T��-�߇�ȩÖ������(���e���[Bkk�".轴#��~,�lo��8��ъ|�Wg��kR�A���[ �5���HaVפyE��fЕ������ժw<��O[�+��e<��(Kj�6��H�@���`{Ìu%H~i�u��s\-��D�#�i
�V�`��QΧc�q�й{��ٽ�_���sDyp�$N$�k#���P�ג��ũ�%�Ӕs�n�H��N�6�`C����~��dZY��!��^�t���'
�����k�9�YA���/�I�n�2|�a�0ö?G�}�ƞi<���"�6�c��"5�F�w��XuLZ��E�%�vP��~\�]rxr�х�pt��HXpi��0�R����'Vp6K�kM,n� �LQl�y�RK3D�<����9%��3�m. �]ٲv��ss��%2}��{�x�����+��|Y�ś�D����^� [^���`dC'�5u�23�-.�?�v�z��,{���TXPd�ja;�б6�C�WV���TepE� &�j��q&L��܊h�'_I����5Y��oD$ qA��1�[�͐�[�cږ�_��8�'E�1`j��u���VZ�5:��\i#��bp0�2q��P��PQ>�c��������}y+�)�h�Zl�"q�zq`���o�����1���I����v �J�e�g_����z��Bu7��Q��?��r���A6܁^���4B��s����ЭOG&�$�A�G��mm�*F�B�8wwV\n�	Y�i���~Y��"��	���695�K�P���pD0s=��JF)���P�+�*��B�y~\!���I(樊$�5��+�� �;�%V:�r�>��1N]M��.���Oˀ�Cw.��I�����ЊYY#���% �ig
-U@�?���n�R�X�1��N��[���I| ��k�;v�2m$C��ѻ�2Vv��@�?Pc8n��l�I+�� �[P�:��9F좜}��
3�W�\���'��$`���_��,�cnx{��ռ�H{�p���WȞh�17�{	��o��c��>/@J�?�l��j�2�a�)��_����SN�O^SEt��tPB��b���I������;?f�Y�k l�{��<̒&�zulH�E��L��eRM8ceyF�%���z��YÔtsMh� ���:�I�^h�	^�`�	�Jn^�(0;����Z� �����ߌ�\�U,����k����O�@�9�T>���6��Z�5�z���К�o]�O�(7m��w�yߜ:���y���G�2���#Zt3��YD�c� V�nݩ�= ���K��9{|�C:2U����
��
(�U�p�f�0��9�:[n�}���f(�p`��7gzџ&�\eЊ���cq��|�s0��,��1������9�_�Q�p�F��piB�-�X�7�P��0�����0���
x�ב���[��g��sf#֔>T-�������g��UB�zg ~���uBE��	��g��gm��.����@ �@�������MA�ݍ��k;g^�]xdS�y~>϶��X^�P0N��oo�ȷ�=��'E��b�F(6⼫R&;s�Ɓ�1\��0:�l��j��mw'f½KZ���>Fu4�'m�7�y���s.|P�Q�4�tClK��İ,�0�o.�i��/Y� ꣃ�ެ�9K=L�j��d�%�<©�҅u'��7�� VV��B�Uw��������A�}.j|+��S�b��YHD�Se���7j4Pk�H����E[�� ��FV�� #�44%bsuݮm�J0/�p=*�/(w�D�E����L�C�W�-��@I���>f�Ŕ �J���rQp�!�	��$�~)u���� {fU +E�Ԧ|�i��!�`�X#مY�=��>;����Z��*? ��Ў�����r�e��Sn
vT��ڎw^g��j�6��s,�r�r�Pz͢��"j�
��K��V�3�>b�\�(��Y���Zޥ=>8���4���$c�p&���)��ò�!�$ FB������4���,�����/���I�Jq$Rk���N�����ؾDl��� �5�p�)�ZD���;
j�r@u�8	ņ^U3
�	��r��?S_v�@Zx��rs1�|y s)���Br�F���t�>�(��s$Un�jB�p<��]r�+�p��iitJ*���0>���}���H�  ��v��x[�_$�����E'j�-&�@�e�-�c�:P$�:�D���(6(��X�h���"׮U���a�E6�j��|Ӆ�"�>Y\�p'F����&������"0���-}�������`�W�h����GȎ׎!@����4��U��XP"�{Y�ڟ��� �"��	D���.��Ѱm۫��	��}8 ���y�R�H�\�u�Y�YS�Tԗ (�xae�Bq4�9�7 � f��r�l�!��A��g:t����!�_S��i{8�5���*����iǭ>�M�:z�(�8��O�</ȹ�n-��3~`y�UN�\K��Cx�)x�J(��_�o q(��Yl\�h1�guu�%�(�|��D�10mE�����TU�Gt �|��?����"���,���"�8,�=���Cmdp��;��� &��~lx��s�&�
ۮ��~uqf$���/A4V̏S��7�F���-�<��-��0P�w�"�Muў��x6���<��͗i�m4��\�کg���l#��E�6 Zqx����"7�Z�߼#���VC�Rq�>�@|�{8k����¿���v�jJr�8cQx����:���ڒ�T#��Z����LuP+h����{-�|D�,6�̓���|��d��8i�E�+E� j�Ff�o��\.8�SH�V^������đ;�|��3�/2O��^�D�@�$C �^�U
qx׍П ���rujw�p���&+k�{ a0� a�����wbzb�x���ot�a�N���ޕ�+!�d0���ik���O�t���������Jfw��{�`G�/���
����r�7�I�6X���El�Л�X�(���>���~�X/Tz��e����{�cB��u�#	�&p۝vN���[ػ��K�2�^���,q���!��
��22K���!PK7"��>�{K=9�ς���=��ʙܧ�j�ut6(m^���0��b��.|�}�o�bN�����z��aP�������pkp���!_xƩ3=cC2�w�+���M�6{^���(��[�#K��6@�62(!�Y�`��-�8�U[/�VsJ0�ǖE�Tǀ**��,5{��)��,E*Շ���	o�.��Q0���{�|�!gW�tg���2���'���p�K3\�e_�3�I�aX�H҂n�O�'��!+pfO\b!��'��N�h�ğ��z�?��|�E� M1Ƽ��!X�����}�?�B���D�� A8ع%���S�2�� ��ք5W�*I��+̍�2I[�k���]��}1��@�bN�C� ���8��r���{�d�Qqyt�3�y���
�ø�"?��Ю����c�"s��m�pj��au� ])��M��͓U��C
���D?RM�ĺm܀����*>���d��>�g�wH�_��(U� ܒ��%�Y��&���p�:��z������Sɵ���Ґ�15���"�Kj_�� x��4tmL�.n��s�W��7Q����o��œdI�3�Z�������^K=�<s�yE1��8H��+3��Z��誌���[	t�l=�Ʋ<{)�\k�A4"�,��E���]}6{�7�p5=�m��%UZ|���Ş�{g61���;���b�ms��y��sf/W���_�B�cp�z0��* �,$C���λ��Q>�@�� b�W0��9�����	*��8�j�.,K���fB\X���kaT�a�X����m*EBxq�,?P�w�ϙb!�M��;���8������f�S����Zj$�?H�'�&�5�vցd��L�0hv�jX�?���؉W{1��<�-���z`���-l�<W��������F���b�u�[�&0���+�������f�B�� |�]��K�c "�b"ھt~�ܭ���@o��"Z�T1Uf�L�)�G!ϔINd�#���v�}����sNV})�/����e�k϶��d�ط� �~�[OBH�O�a����*6�lj}Kp9�"��Y�l;i�X�}��4g���bqށj���W��Ɇ3,4ϥtqN� �˻��$��
P��_�'�i��o!UAh��l^iM�m��%�"�_]��S�U3��5[�X��{��� e�H��ґ��
�`�՚*-@�yߝ�ei@^�N�Y����K7�<'�ἒv�|�\'�l���uXF��Q�e]�˒�|n�Ǧ��t.�%	��5J�s%�(�I���&��'�������"���uH�Or�`M����_�o��b�N�_'�zLx�(T�"�0�P���N
��� PU���D��P^�;sz���P�&�
M�8+���\˿����O�ϡ�C��MQ������ΒR���7Ɔ�������Jn#�Rd�+�-���=f��r�-�5�p^�����O9t�J�R1g�b<�;���H{`mT����,W�<W��J�ぷ�N���/^��7���ǝ���5�U�A�d0*6ok��v�W_�)�]|�犚Y������=���b�t��e.�iYE�Fd�|���w��-�R�ۤB�J�X���&�(��Ix`*�")Kn�TVX~y�y��� �Q���cqVEYЬ0��+9w�~~����A���R^G����g+���盛�ɨ���-|\z+ל�= �ɩ�4H���|DSj3{�3�U4{���,U�9uۀ��mc�Q�8u|	���3�Fw��T�b0R8u�U�_}���*<���v�E�Ý�`���h��,��z��B*�I1ܘ�3[!3�6�M���q!��d�.�{C�9/_Qӓ�`|�SߐI�rZ�F��?�ȥZ`L��� -���bbG��f,Z끐L�qV��Ǿ��g�n���� �xއ4���2�5bn �>��3���c]�����e�B}K�`;�	��Z
��h\j�����4�ẳ=gⒸ��g'���G��g<
'��'Ey �7�c�#uw�0�Yo�g�5�o���}Y�9L+��Mh�vm��#7���XA8 E�M��0�*�~����쉳�р�5���ўa#=���PYӗ� ���N�=���U�Ր����\LG�u��.��hiV��5 R��p�u�U����N�q��l1������x?��R'�65�A�)����V%�� VP�ރfqf�k0�͖�8�[e�CO��{���n�`^����ŋ����5;ۋi~b��§=O�s��M^W�Tʊ=2��͙�h�+&�]�3IA�o³�[���<�c��� �zd��9 ���]I�ݻ�u���wP�e�����/�ε~4�,-)��\�F)w�s����̉Ó��j��!VXU<�$z��t_V[�Q��!��c��k_V�/@�Es|���R\�g����ɰ@@w��wH���?�����b�B���z�m;�M�cBT�~�O������vR_$쪙���cl.���D�*�^�ߛxM��jͧf ���]	TSԻ�Cֆd�M8y�T����~z�c=�լA͡X�RHȜ�=o�=m�?��y���s��B���RRߗ
�l�=ή	�գ���-(�!�s�ɐ�a1�s�d��R��?_@�<R��H�瘙��,�����z/c�g��Z��f"��K�g�>�Q��E�>�C%m�ZbQ�.���<u1͠���ms��MVY��55�0�x��LAa�oz����f;K��P.LgCV!���?2#�)8��ч�v�$�
�{a��{���g�h��N��߈��t�1^�&�����K�y��y
��g ����K]�<��N��E�;~p���s[LW��M`IEj�o�ԁ��~{� ^��N�۠f_֏a�8����.�n=��wX�+
r���L�v�-����kʙ��C<ϰZ�g58����\"�{��S�w����k�DQbR) ��cB�L�\-q�07�Z�}	�w�e؇�˰
�)^��oB�24h���#��:���~?XZ�6�[�����cQ#���L��D=�(�@]�;�JB^p�?Ox�Ud��!��A�����^�㓶�ȫq�l�s.���V�`�?�� �����EWA�T�{��8�HiH�;�y��ߐ�@�=�&~�R%���2U��fC��=IY���y��T}e\T���E��"ҡ�
� 
�J��JIKw�H7H��t����t3t�0�4C���}����;'�^{��Ͻ3�H��t��OwǵLT9"��Xd����9��Aqf;_fF�1{���L,Z��ن�e�V�f��Z{��<�F5�@	�n�R��؟�	4{���q'(-��U�{���w� Y۶zf����s-��U����2)����`[ \�^��3ufo�ҿ9�HKUr5f�=�Y���6�XiI�.�nIu*pT�g���j�y��`O�a����0���:'���{��*��Nu|���d�������S�Dg�6I�1O���E�nu#W3z<Au��{X&�Z� ]�8���B�^i��Du��Ň�JY�*G��`E�6�'�=-��̀���/�tqޱ�O��{I��oc[��S���~yv{��s���jx�=O	��d��`��11q�D�.}����ͧ���	`���w�D���o;�tV6�{K�#�_�X&@t&������¯/٫O�A����"N"�ľ�X�j||H�oj5���_��m�G�YOL��[z��=��=�}�n�l�U�9�����gͰ�[<D'����l��Ь�׬O�='Fq���"�+Zrᗨ�Կ:�0n�z�UY�$,�$A�C�cgĐښ���L�/��\��_6�=�z>d٫��w޿,��8k��G���Puc��I|yK�{e�L�_�8�Je�3���e%0c�'��/kŶ
�U�}�=�EĮ]�����nw������6�CA�	jh�9{�V�?L�I][��fz���&�M3�ƅ��6����I�eF�<�k��5����F�0߁��'��⿬�j�?R^Q�?��Engf%�M\������WT�woS��=��>Ul� �啧����Ox ��
�z\�K��0/�8���u�q�˃գp,Տw��dG��S��6��oSAIj{p����G���ŲV<|˙.����؎�Պ.g@����,P�O8����?�\���}}G��3������A����� )�Èf��(f�|t����Ѫ� �C��z���y��A��=7���n�\�^**����&�Xu �)�f}�:�|�Z�-�z�#�3M��Β��"k�VbvR��e�[�[��󛝥�	�M`���������g��}�n�SԮ�>���8[�gI!v�{��A]8���rDu��>ǿ���9q9,Q�������f�$�C/�U-!�������6���V��A𺌢�́�5�&�؈[�Zc���rtM���T����n�T�&\��	9�=[_����	@��L�ҳ�JV�i�������@|���񅯔��:= ����A_�Or�q�
���	������@�Z��u�&�gT0L��AuҢ���U]y���3�;_eU�i�����Z�:����+�cq-����2uN�v^�`I�{��A�3AR�}"7d�60�H��w�5��i5h�t��]`|�ف�����L�:~��VS>�=��e�^A��gu��y�&hL��YO��A�)���K�|x:�b��@-��ô��8p�p/�UD�	�oW��P�Z6�ʵM5B�8�}�
��uD��Eϊa֖�_��3dtl-�fɗ\�j�>pȲ�o�1s^1�b�
�i>�^0�~T��]aKD�}�k���hN�H�?�����TU��$��*g=,�Զ��`���=�z,�@!��H�S��#.m ��~�^[ͧ�[����J���{�Jm�����a�U�|�`�Gw�����|#4�ز�:"Fk�����]ѓ�/���ѧ堝�����т�c�;ίs���W�����-)H�S׿>�u�������D�IS��>�EJ>2�~�*� a��������#�)�r"z�/�0;��ۚW�h8�m����.�>��v��M�Q1�;G�z�4΀y�9�Ïd'"��R�-������v*��=zv�'���L�t�wwS�&8<�2�]A�t��1D׸<�J4/Ɲ��C�Pz�kĘ�9��m�838ht�F6Sp�#�� ���>Q����56a���g�pnnI��u��V��nIAw��JZ����}!#�ݕ�-	���S~�Bsp���R~������� �����N�o�f����i|D�Vr���M���j��o�qV�P��0��,�Ho&N��u��ȅW>�J�rV�8�����K,7��L�D'	��$i��ߨ\�8y�RJ�;�U��+����Ƴ܁8��g��u�I;
n��]ĸ�q��Scky=S=ɸf����]���c<�eN�߼�[LF�����q|-*���|$S�,y��%Ԩ��X��K�ۢ�wcŽ��[K��ݣ�}*_¨\��(�<�Aq�	��T�tZ��\��78���n31��v}}5�'~����z�����N6�/���%�{ߤ��}ZB�K���fsiR�?��U#$+£2���8�ʝ��(�WP�L��!�,��-6��B��lr��	4	�	K�"m��:�fK2�� �ܩT���\������Bn
�;�]\�|X����;��1ƧɜQ��#t�]яª4����#�yf$�	�Q۬M�8(?�z �-�^�Uc�ht}�_~��V��>d�L�|Oor&JNz�е�sb\q�:���E͙�v���#���n!��u�S��
�}�3^���;��v��I���t����+�Dv������j��>X�jܔ����3tv"p���bp������΄���r�Q�J���@�'%R�&�jSp���U�,�_��/�{���9�'>to߹�<��N*�m�8J�9�Q��Dr���׫���g�!����
��g��^Րx�Y?+)�1��Φn�B�~1��I�֨��%b�6~�dﳭ�|���6m���L��d��"u*�?�ܻd!�1l��[�����~�{��k����욃PL>�\m�l�C�軕^���<��]��F�8Rk��WA֨d�涡�n�oJ���ֹ	��o�/�݈t�O1Cb�A- ]�Ep'S1<� �k?O����v\�{v4w��ONd8ҿ����o�
ADp�@�H��q~a/�+������|���ߍ�E?4�`s�뉣Y媭sx�0x��oO���֍D�;N��c�e�n�bլX)��KuJ�W��I��ӽxb]���v�NJ��Y��G�5�r|�w�{�v�	�$ܒ���p���̭��;���28E}���j|6|���[��S7�¢��w3,fR���A
����v	۽/�Ȭ{k��:&�э�}��ߴcdy̓�lO�'��y�� ��,R�lq������T�Ǥ�ʝѴ]K�z�Ӛ������I�;q����?��(y�>I����]$:eW�eP.=j'�����~�}�j�,E�D�AR4��p���'i$�� ��9�T�w�EI���G���T��w�� BǦ��U��
�F�zQe��}_��{�yW�:+��I��K3��hcwaҍ�?�$�n�3�J��5�ŷ����D5�P���Z���d�y���ᢟ����l`1jt ���mt�,S�����v߼�"���O�П�]~�5,C�KV����EB�y���1�s�Pseh=BܻnH�9���&
��j%RD�<���3��̥(��?�P��hv�!�W��C�]�������Hi:poi�f~�9uMY���th���7�h/mu�%g�Z�����T#	�7���\ �3�+͟0"�q�������y�(�ݗ"����MEb��^�JJ�VH|����9[U���n��#n����23N�C��=p�Om��cAe5x�X
�V.��A�>J�B�l���_�	Hzч�{"<�� h��/BĈ
�u]y�9
�#�jZ)�u���]��uAa�֧Gq��.g/ڳwH��-�#0u�<T�݂C7�^y��n����K����(Yd����n6�&��_W��ep�����ބ5�2%IB��lfE��d��_&������h$��LV����
���Z�	�������:��HbX��G?��?}���ۤ����sv_���}���*I��p�IMF klbG�4����[����ټ�@W��|��:_��)룶��Z����a|�OxԘ���ї�B�N�ry�!o��r�$�%J�o�Ϗ>�=u}s�3�E��'��F7*+���篞���a�ebNЫXQ��O
Ϡ1�ob�vݹ>�-v�C��}3�%Ue�/��Ѓ�7�*��߃��E�ޥ��c�c&I�~Jd��:�Cvo�E����މ<�.�U
����{��ua\�}Zf�����Ԡk�<�Z���P-8Z�\(|�����O�������w[h����@�}���lk����ݭm��w��7��m��A���pCt�o��0�zY@8�GMx�+���yͪox�@	4M��j��黓x���_�%��H��w���c��jYI�'�E��$�@x�@���w�J�}�E�BK�?�)���G�Q�'�b���%�<5?�|*J�Z���Gw���"?<����V�=��/�S��{r"��йbf�G<��&��I*��u�b*��S��$�wH�	GI޲qw�����A\�Y��8�L�ٸ���5�2��o�C��3�1�H���o�
a$�$�+��&�(�`M#m�/ӡ�T��j�v�4���	�����gl`lΧ��8!2�=�:�d N������~�Fr�V,�.L�.bY[�ǩWK{�U2#K� �u��Ԭ�S�{�|��&fը���[��%�LF�&��)�/Z�H ��N��+��#��k�ya'g�Nj'���H�I�l%�r�2��}]ӑijxt�z3�	���k���ۥ�?����\� <jY<hV�5�؛}����D��dA{�4-��Iy	����L��ت�����s'��s�������2I��Bd ��9�K��xuWF��ָA?N_[�S��D�G8��t��6������)��`��;^��\�D\�9��"�t�����L���W�T�L���t�'�t6�B�It0�Bv���G�nq�Z������#i��`6��(A����Q��3=�ãl�`q�v�J� ���?��/�)5��UO�Bid|9�?��9��-��v1RO�[�"��_fv��BY@���@S�I��>5�Ӹ]2]���y`��DV���QU�3M5=�����Q��o�B�?&�� ~%�5&Z�!�t��?���X��.r��� �_�EdH:{O�Z�{�h�&�da����'����I7lUy;
�?����y/D��l��j&V輶��p�ܻ�۷�
L�2*wI:�_�l��(�n~�-�I��'�.���J��r��7���P�r�f�iRO�EK���
g2�խ\�;)Adh�٦�1�a�QJ�\n3��(���jf(B�<Z��y�������|<̋����=�ί����gۋ~ܱ$���8�]�!.�i��h��I�fu]��'�K\s˗��V I�N��8*^�S��q��� �у��p�V��/���o�y��w���I��M(qH9��� vT.��*�듲�8̖;Þ��qV��Kl��J�m̅�J(UzҚ.�'fe�����,\aLb�����5�ԍ��;�u_z��N�t��WV��f�����4P�ͩ 5�1�>"�{yZ�#tF��c*��xo�o���cF��Q��s;D��c�9���).��h`�p���\�D:�{b'�8�2'�FñȖ�3cV;d9ٱ�y��1$F�a��|�mJ-c�H�#��e�(G裯.̉5��a\?�,�Z  �'k���;\[%��h"�;/�͇��f��C�t�v�Lbj��� �����I��07����������
vM<�?��_���J$x�<���h+��A�9���Q�g �9^O���=���Y�|��t qB�>��v/9N�o�0}e�2���}�\k+++��e �B%���u|���Y�|�f�z�3�Q�4�Ө��Qe8��oN/V�y�d�4.���-��&��s���7~�W<F�U
ð���ny�Z����u�s<Yl�ˎW�Tk����2����Av9%����v�l�|S0z����$i���Ev"��BW��A�Nɫ����
w�_b� ��E7!vJx<]�L�u�wo���BtYR����kZ�0[�먂�11�m�H��c�4M����oԯ�E"w�!<|�9��k}^�cN�",j|���|�_&A���}��ߎozlG׺�<k e�g�U��@v��ǋtu^ښ6>�����*�Ά�U�\/��h5�W�Wx����'%�l��q,;��ק���І8�ʧ̷��	<�? �����A.������,�1����v�B�hgC?�wi�P�3�~P�y�xS�=#�+#"����߰�P��m����FQ�$�HaAx����ͣ��|&p��I/���1y	V"��	�BM�ub����~l��4��_�`�c��Qe�x�ȟH_��F�^<�u΁ց�(���*>�P�[Hjňm)-�_z߹�S��.4Mk�q����:��A��<lj �%,"�B\	.���3�_��ܸ�ԏ=��o��6mq�L���!��'$��T���ĵ�5(�}�&s�+@�t6������{z/
�}�I^�
D.�A>�aj�xGUJ�v.ey�b��èAFғ�\D��^��hC����{�'��T�ɠ���Z�_~�Px3�2�7��_y�,'���浳 ����Q��4�h�uUͫ�E0��`����e?��P�'���vL��v�0�0�8 )�bW�^z�/��s��pո*���b�ar��˯�?��C�J}�j��u��x'Z��@�ZZ�(d�dL)<�7� !����sJ%,�8�6OY����l1&��?0},��,�r[����q_uS�_����S�^����i)e��N����փ��0�W�T�`����zRO��v,�q��x`b�<K�\�r��U����)p��ܖ��j�*<L��_0�����2��v�B��3����zg��t#���)P��@��;C��s�~dW�x��Y#��J[�O
��5��"&�eV�)=8��ڧ�5����jbZg� ���������kD\̸����ڬ��ԩr.���q \�]���oc���&2@����ȶ���;��A%-�з Pxͳ{�?ʽ��Ռ��#��trk����_|�h�@К}>_���~��3ZǙ�M(RG�|�`~Ъ�Up�1~Ȣ�S�sK�W���%,:х�X��L�qfj"k(m���}�;G�O=W���h�\!T�q�ŏ�$s�G��r��P��V��/��V��u�����qJ��)��4��mY��)]��?j9��I�,�&�*ssF��_��m�1�Lqi~y`��@&�*L@&��'1�魹U RF���5X��������
+��,h�fzG��B�C�5���G�%��G9b�7�F�4��b��S�/�J}��]��J`�V(]I.*� {	�~-�!�.�s q����˰L<�SORt��B`�׶ lH�٤���3b�m���ٙ^)ad����8e�c5���u��0$��PaGl�����Yi�P�F��BS3�������]�����a[��������e��!�=Ѐ����&�*�9��ywD�>� �y���>��zn/�ݢXk�� �O��(\��<����
Lf�?m���2����[�#�=hE��fӾ����겂����:nUt��W�9RCt�ʟ=��ώt��oU5��&j��Ko %�g�X��r�����Yq�M�i�OWӕ��D ?m�����eg*�����(J��'1�j��U�6
u���i�>���qeiY�]�,�nX�Il�H��{���|,��n�f��ʭ�te��J9��OG��ڱX�^dV<�q%.��Ӫ6���fE["�˝.\��Jf��d����p��p�����KI�
ܗO]��rS�}r���M{�����C�oU������[>M�;�J��B�N]�A}{^ ˊь�Ens!Vh��K�4t/��K�+���Kr��
q!>xi��yD�ȗ����v�D�K�������Ж��=��_}��lΥ��&�W�L��~��]aYY�P�ϡNk�A(�+I���>c���z�]��+�B����'�V�9�57��v�F�]����򩦕���v�����O�g�P������X�itKt˯l]���w��-�}
�����q )B��D�!���Q��Q�T�,�z���W�����L�yel�)�q�$ߌw9�KǨ�E(�)~��@���P�0����ޣ�{�#��D�M�����E�v��jg�+��N�㼐>l� 9��R`��\��Br}�XЕ���\8�D��������x�@,o?��� �S���e[�w���i�rn�[�?�4y���S曪��޲B�����q^����V�ZT�3胛�tY����)Y[��eit�1?�=�OO��	����D}��Sڈ��k�W��I�z��j�x�&¹*����⾉ڊg�3/Elxރ�� ����� ����nB��g_�����+b&���d�W�^����p����%i�O:���i7�Gة�v���6��r�ˈ���`@���6�^{�qqZ���c���(�X�'s�,����<�b0B��EE/�����_��pob �����ϥ�4�-�B\~po}���z����m���Lq��7�����9b�Α2!��U�nR�]�qH�C��
��p��y�)g��<�����GZ�f��Յ�m�b���r����gj����QU@�,�&�f���H�<�OVBER��y<��d�~0�D�"���Է�Q �p�i�3�vS/�zX��wF��@ڈ���=P�洑��K���U�a侫RY`���
Z$�}IQ�4���|#b��^� �	��8�>R�'� �Q}��y!�u0�[@5? Y���y�<��WL�dSi�H��Tkc�rH��Zi�r�6�N����SMU��3������3�՝��^����x�ݷ�Y�D�$�g�;[�|�r��^3X;�A<ȈN^�M6��+D ŰSV�;i�_�U('�@���7&<���v��OeD7J�:���Y/�@�g��̑+N�X��>V��n��ju�F>Hz�0Ģ�����+���.�v,D6͌r8�v@?mc����6 �T�#R�'r�Z��	��	/M�Ęu`w���
�:���2:�����U5o� ��n4-��T��%�>��fh+Kؕe����J��ի7��3�R���g}� ��K��CD-����	�� �.l>ӕ(ܻ*t?0��4�r��3t�\3�Y9Z���ޓY#@�Q/�N帴*o͍�J#S+[!Q̤��d��>t��[�q�/t���{l��C�Z"y9�!F��N�.�����摃�	(d���Ξ"�u�D��ƗUN������N{�����_ܗ��5[l����N�^���:EM�Vse���ꖈ���bn&,=DH�#`�v~�/�(�z�!��[/�Ҡ�ӈ��$@�Iw��kdB@P���D0���[7p���|~��=t��~!%�Up׿�k�TkZ%Bd�[l&��>��$�!���pJ冁|��^~�<����7�d���[������g��Q!,I��b�2��)YC�i�k��+mV���I�wa$(ԍ�M�D���\��}���Y�� ��v�/KI(fe������u�_~�m���t�>ȴ����F��xq�}��$�L��S�:��]<��N�zVp�M=�������LnW)�(���]
��Y9z����u�����8��8ҁ��}���*��<�}�V��~�۶0)��B9�@��~� �A����]��,�v��j �����*��#F��Cx�W ����p&��Aq�z���|���<�ޡ"�g) 0���<D�'u�}b�si�z�W�|�������"����;��R$Vt���O� *���J�.}�N�r�m�TSo�������L=���8(���7��ys�a�l�n,�'1��@�����_��L��;���OpP}���h�A��1$s�3�o/��P��61T��B��ԓC4�����o2K��<AS-�a���d]��-b��*}��8*��V�
�́��V���OTHMo�0AA��L�SG����*��^֤������"��p�1]I침���jf��g3h#L���6��E(�h�1y>���ѡߙ%F1%���Ӄ�'Ӻ�i��!1X	� *��͸�,]=~�:p�A�g��+�\Ic����d�[/�s�7�\yk�Q ����[�h�L1.R,,�SC��-L���3^L0�Cf�}��3��[�E��S8=dWSx��0��=#��*��J�?���?�[OJ��ܭg��Ѭ�^d���s�x<u���(犡�z{�'�J�K��{�7
v�I-o�����_�9 \5ÝO�3�2�ش�'W���U~;d� �(�I3�B�d�Fl�"���/C���_q��;}���@"n�^Z?��@���2��BC���س_?QbV�������yb�����35����>}���3rY���Db�� �W%���N���~�K��X��AK�/H�\=�Kl5�Ĕ�m����?�LKhY*���|��d�1Y��H�k��w?��̤�:�|���ֽ�t3M���[}O�Y� 
K�f���5A��Ĵ%�4O��M�������3��;����Cs��e�
\�뱈+���=N ��h*˔pHW�$�A���̩����� �O�_�zO�B�����[zU�~��ul:ލ�s���y��Q�W�P˯�2-�ݬqG�Gvp��ᓘ���-�W�ֲ��7������s=�f�y1�E�w^�Hy`1ů�`��k �Z�K���K���/I��m�+�˥E5j���:��h
ÿ̜�`#ɱ_t��N�s��{k��JNZk��fB>O��c��H��I�qUf���C��T4��B��]=�h?5>��w)�q�/���t�������|z̹����l�$�Y8g7��c��ؒ�<�����%+*�a��e�bT�;�ڍ���Y��V�<����b�X(Dx���(Cn����'�)���M����z� ��S�A~�XӒ5>��W����)��L���;⋞�z}��WC�u���R�,�n�ӃOuhǦ2�DP��D�nB��g�?C�9J����۸H��z�A��������A>W�\�U���΁�E�<V5�6ޏ̢��	���f����UH�ؒ��o���D�;c�5*�16��ȃ�"0�d�^/��>8~���� mL�-`��;sK.T���$U)����T��}�=����!7�{=�r��Ռ�)Zʪs��^	�h�L�^j�_ZU��3�ZvFz�=��(0k�ȁV`	O}A�,mi"��cL0v�����م?z�hg�K5��������	�V�������-#��xJyTvy�y��J���d
.@��EQ�~�b��n	�N�&'�շ�C��рx�8���?\^
97/V&��g2�����.?0rǺ7�PJw�?_��tY'6��mb�qk��T��ޗ��p�?L3ҙ��C_��`)�P�#�d5�q~�؉ <n:oxy�b�Q�̡�,�'+���5����]�If���p���K���M�ƨ�̒v�P�3�b0�X�ਐeZ���w�VT�,<�j�K�q;pl!�E�����qꖲ�;|������!z�+.@�����c	N�؉Q֦��h~'�4v8����*�}�^�B�_����[�c��#��	BWy�
�[h��J���~7�v'�U�rq�E�1wz�L�K� J����<����h͝pT��V/��k|��g&���9;��K@�0�>EFD�����غՊ�~q��<�K�wh�O��w�7<�G��
Y�Xnf�{x�sSh�g��l;6��kk@��vz�u�c������2�C�c���������{c.���3�~҉P�����ݧ�4�q���.tą|,����ÁecD�E�l}8b��>��2�A]�p����\�QT��N:����Z����E�ŽV Ŧ+4�|��u�H��{����Ώg�R�Ip��M'L-�3�1Z��Dn�&��g�Q�M7�����%���u[M�R˘"+��^ ��Z�o����C��9|�Pq�r�����j���O����VP��L�+�lg��l�z�X=������m^�]���Ѳ��Ǣ��e��ezV����ؑI��� �⪬Q>h4�hI���Ҿ���\R[GZ팀��&���W��g|����yhX��p�e\�.���oD�}� X��`xl����e�{I��Wr�V��^	Ka�ʯ��/8G���`y������*��~�Y�פasK��Ss#i���\��ٞ��Ű+���C*�y�S#S�K$-|�VG*:A�ߝ)&3��q�(�b�ghfINy��$iK6Q\[> �*��u��q���ĸ
[��
-�?�nٷ�{R~��{���b�)P0�R�����Nn�^I��i0��QRB6ERsw��ML�8��������P�^&�����g�M�;�'��#GP@s�f�J�~����ܣ��Qܯ�r�O�΢���y�W��`�]e1�D�������uu�h�� ������V�
_ �Ң�Pyv5rL�O�23��3��v��C��%�u�g\1z�4(�v�N9��悥��٤�q��>�xQ��Rb_�UJ���#�A�;�)���7�+:D#����"��@�ã��rJ�%����l��2�8�-F�Q�z���Jq�J�ތ��h�R�`8f��}U��SOvw{d�C,J$<uӰ%Z:�NB�!P�5���&&�<$��V6V�`3Qr�A�砝q�">; ���VȨ�/��N�?��\�s,[0�	��v�L��٭t���l�=�����N��*��1��x)<���a��$�Pj�a���w�Z~�ï�kF�̨vd`@%\�> o0���
��Xk}H�HO�e�(A�,6j�;�P.���.�קZAQ��j���=��u�R��S<SU'����V!G?�k0����`	�5��TeQ��t��Dy@�<��O5��qՅ�ҁH\(���t[�q��ǐ:h>M��F.��O�o�]�!�|�擷��Dy�>UM͚�X]}��c�%�:XN.�:s���~��>$Fm�=���X[�����@�����$��eJ*"g�v�<���x�=]Б�����6MG�	=��#��'PCl��#��z��۹�d���z?g��I�˫�9ț3#w���t��zϔ6^�g�re�=jhI#ڥ�-)~ �e��8Q��u{j�-I���o<@���|J���t��x�>bY�xt�:p���ܢMѻ"��r�'�\������l���UD/c������I�Я�,GH<��!�ثa6	��&^[��� ����)|��
����H��@�xb��V������ɽ'��7H>m���WDj��#b,cR<�r�˺<q5$��J(�l��kC|F7m���U�̿�W�)]����B-'~�@�-�����-j�e���?��]� �mw���l�`�a�u`w�7r���+�N&$�dp��x��"{�0V�E��f�x=�����^C�+�g�8�:AÝ}s��Æ�,1����:�ڊ�)��������+�y�6l9[9������*:�	"�6Յ������������@D�sp8P���"��� w#�ϙx��R�͜K������R.����U�7}����RzڰM��ە��{����D<�^]�C�<.>>ƅ���Q± �V����Q����ż��(�z~j�o[��2�3�a�fK-5{�zd�
��G�x�%�]�����TP�+��Wlc./p����5��Z��H� ��b���n���=�lf�~�v�/g�S���4�^\X�:��r�cހ��>}S��k�kwe�oZ����^4�{����!B�k��l����S�c&���x�0���
�c�U.o��t��Eh��"hF�p!H��,Ѻ�b�m��1b�	��03�ֆ�����'b/��>/�j(�O�y�ۜ ��%=�h�i|�����٩�h��%����)����y�V�>|b9՟��+�ߑդh�jDm�������*~�����G�̭�w��U-$-�'"����P�-�r�
�Lf^g�X���|�p�Uic{�\��	꾝�þ��BA�4@�=�&+��pԕkԸ�d�ص�H��� ��#:g'�/����KR��+���?�k��ɞ��Ƃ0�	N�o�>��+���w߳Fa���С���e��Q�9)������*�}\�%��gL�z��o!��߳ x�y H�0��S7�;��,�
^s�.�GM*ϗ���G3w��I)���1�!_��v���v�@��T��� 9)�w[���:�{>n^���VW�߿��j��)y�Vc.���`Po�-�M9e[ԝ�)b5
����.,R�,�D�E��*�q�W�����Դ,x��F���~'=�x;t�#��r/Éϙ6r�,�Gϥ/�E#^ ��nF���p��!�Di��W� ��7o�2�l��1~���0���aඨpF����� Y�VjٖX�KO��<W��#0�M�����G8���ء�RD
+��	Vh�WZ
r���OFs?��M�D{ͱ�y��G�5j���$�[���/g�����h��dd�Z`/#S·�	�f?�����s
���w���ͷJ����m��?��;�i{s���A�5�7�+V���;�1��y{H~ȩ�Y� V����+�9��6��39�N_�-P���7���bG�M�d	!�'<��{��+�,�Ͻ�����6��F�6/�@lg' ��^�)��Q[A*�Rm2*�3�V�2n�d�4�����]�{!��!���èi���bG��#[�g�ӕȔ�)S\�}?� j�	����}�뢆|.e,����4B2.�׉��~e�_��0����7�I�|�\������Du�R�Ӓ
�H�óA-8��+��y)I�8뇴���;Z<�#����c���Cr�����;=�y��^s���bac�[�6�VD�>�kx4^ۏ2��y;��z���Qy>D���t��hO�nVT����fF	
�ҹ�����m�ȊDu8�
�m���^J��9�/�⬠�,Ϟ����H䕕������Spsa0Wi+Bߝ�#-˫���䗏!(Ԅ�#��2�l�`x�Ǉ�Q�zq�o�ٟ_���}�ls]&|L��c�#��d}�:�{Z�z/ ���w�^CY.�ڱ�2-O»vC��Y�?�	���|�o�M����}w�H�`��^c�dt�7@�2�ȧ0�kp�j��A����5m��}6���ߟs�A+��ʗn�oI�9�vY�����n��������*m9.]d�X�Kd��G채HF�#U��VGG��n�z��&իD?��à��}`�(���6u9���`��M6�e��$9;���k�?�{���sb��
�e;:ei�e��D۪[k��`q����+�/	��(�*5U�t�����H�o�AY��,�d���[�/@��\�.�k���Ck7($�ٸS\���������.!�A��ϟ���U�ma_ pi�f�7{Ԝ.�l�s˫5�6f�N�!6Y�������6�w�)㐟�gZߟ�!�m.��.&ٿF���$�\��8��b=�x~���׃��s�&	�"Ac��JWz�h����"���V�J��KЈ��|��R���<�Z�ԁ�x:�¨M�Mk�g���iYiy�����9���Q����(ө�0�z8��&��1��dx0E�������%5m���R��VW�c,a�����kjk��8����ad��=����h�N�f�/���q_=�~N���C��7���!������=+21�w�ʈ���r��_�w�%0�j3&I�p�C�e ,k��-c�A���Fߋ<� Mh��y��(�\��H8�o�$�ld^���Xw���E�dkXU��S����Bt�"�Xׇ��Ƃ�ˉX�^u�Ҍ��U*�yOa�7�r	�z��SGY.t_['>�~_kE��j�V7j�Z�bƚ�����E���������T���)*]�ގiT6�a>UVO�s�95.@�p�}#�]��L�_!bWȝ���r�m>�p�}B%�[��-|��k�]�*E�6�ƨ1�R�f����E��z3B�>yg�*_�1l3)�;��v}�ӻ�k��P��gkӦ�K��0/��(^�u�kY_E��rD��و֦Zc��nC�}g�m�# ��8P����^#�[�|�u$
�W�i��>���ZN�8�K�ڧQML�7W���ة9ݞg��;���9dd�T���sn��KϘ'Y3U[[Y���TK�hN}O��c��>�t$:�|���}�\c��ȥ}	F�CZ��3��«_��v���.pj�A�(``�[�#�_M�>����r��1�F�k�N1�X?pc:}��xiI�P� �Kq�r����˂f�Պ�Gޕ0ٰ|�o�~��8Q�o��]K|��ɐ�W��������զݍX9օ�{?&|�����W(��
�)�-����@�gG��+kO���H����Y����u�5�ʐ<;�ţA?P��CCS���d�%a�5z�:,���+v�8Ԧ2�3�YYΈf�s��R]I�b\FXq��B���0"hPϡ�`Ёi�$^~CQ@�Q��N�y~{�������r�t���(>�2rJV���j"%�-)2U�uvL���x=�j)��?�z:]-F^��$�'���,��'56>~vS.:Qk�_��G����x�LA��q��>�n^R/�yBeO��p��̦��_��}��4�jq4�e`2��;�;�xS9����J!��:�������'�������W�)���� �γ:�_|\�{A2H|@�5�v��lb�`��͚�g9����b8���wv�%.	н��ʛ��:aK����d�N�I�9{���!(��j��gJ�H:H��$6�f�.ҽ|kx�[���@ϺY�Z_?ƆɁ�ة�5A�Q�k���jL�(C���ţ�
�rJ�<�H��Ȕ*IGO�ؐH5ZBE�0��X1S��7p�A'�}je�wƜZ_Ѳ}籠����; ��z}*����7l�Nk
���N��QM���||-k�^l��0BMj���� �3U����Y����+���٭���BB�r=��Iw_��t�<Ł��fP��Q,E;�~Wv].����������r�����ܛ���3��-�r�!UQ��l]�[f(�_7ݱ��k��eDG�)i��
�p��B��ނ���M���p#�4zo��	m�r���au���;J�P�MЀ��=�6"���8��'������~ ^�x��F8�4�.��Ϥ�g6�q�wCE�b�3ծ�4���m`Qm]{��n��C@��n�i�	i����t	HHHHww����~��0>rf��z׻���ٺ����/����z��� R��wn f�C�C���?Cv;= 8iXV�t���z��wi&�+���ue\�]��)*o���Q��j	�����kt��oDP��ޮ 4#�.��ۏuT4�N<n�.d/�1��a�;D�	�m����:4*����_i$=ߟ����k�	���ɡm��9$�HV�9�!h���b��Y&�2�s�k���|�6�\�㰽������2C,���^���D�����d�i܍Ⱒ���nam�������' �_�!�t��3$����W�w'a)䢇�B��ٌ'��7�r+��Ҟ҆?'5����S��kd}٪�;Zr�;���˳3���LS��~�7�l�����$;c���h3]%�à\9�U%.�};�b�=Q#���@��i&n��Z�/�֠�ܸ�;u!*�%�"��l�=���.�� �ט'7�SV+��g�(6��U?ņۋ �o����a)���gHݵ�@[+5�*�B� �WN�ڶŮ�Yj�bz���ɐ�&o�����4[��84�e�V��6V��ʐ<����.Y���k�2I� �(%�q&K5��{�nb�k_O7�^���A0y��7���k!~l��M�A
�]�ݯ��6HU�W�b=Ԛ��Hk��Ø��2�z�n�'i~�m�#~����9(�%v�h�`,E�M9��C-1�_����Q�;R��-)�{z?>�r�ܼl;~����qf��
Ҹs9U�52�/t<��Ap��f�O�_���<��U�cL'Z��K\A��HalB��JO�V%C,
�7g��( �r
띻���\r�w��}3.p��W�Z�lhlp|V2��P���R���Ͷ}v=[�ĸ�����x�ї�~�v\>n�4�v�!���;�
�c��vs=���l6�N�f���7��x� ��w0
��[�^���|�(& �U��V����xms�^�O��<#���<�r���io���p����=*�۹����PX2�)�Vf"�}���d��O����W�ֶ=�#Fû� �[5V���U��X��^d@9���������l�dm���Q,7�P�l�PJ��/�ˑـ|�/�&ȼ�Q����y�^�����f�g&+����R���X� �*p!nZ��k.Ǖ�s͗�w�G\_6��F�5���ٱ��#�M~@�x��	b	�-����$�|oӎ~
�������<�LFE�p�V9n.�o:����Ѽ)Y���nw9ˬ�4�3�ex����������\��G*�M:6�:��mY,O�05n;���iv�*�Dʷ�R[���n`��I��t��`��2��s���:�k��r3R�Z\�T�07&��]ey(:�z�r���ت�*�u$���cO�I.N��᛾N�����x���E�<�"ϣ�7�	�͟E4g�؛�-F:�sQ���n<|6w�d���D�f���ttJ�Z��{D����k=,��k2�K��ϟ���G-�|�ݯ��X��@�T�w.�6�#��<��pt�ԫ��
	wģj���Nυ��`��h��	�����'6:��ꋝ�9�(c�l-Y� �v
�b��sE),��x4oȒ��?l�j{�/��5�;?�lv�e{`���OG�V�L*������H-Y"m�p�]��֤s8��g��`ǀ��˓w��FK����F��_�EҒyA��B���I�_���,)�W8��11�tdDDb&Zt�c�l�b�]+3Ƴ��9��/�,	�M�6���4j��]���$J��-�P��f����;5u'�m��4� oh�ţ��1�,/s�Л�L�7��C��L��_'*!��������r\�z0�XDDR`Hc����ʸ��><�)�E�e�k$�3V6(I��:��� L:�xx�_6�-xs��j��4W[+��+�n������d=-�L����`!�k������J�^�o���b��Z5P�O�c���';3=H"���_��u܊[8�Ҋ��eI�)M���n(v�P���w�NW?x(ƛ�8^MbbJ���S�А���#��z�s=��]�����������Eefp�,�o{c}��1��X��oZ�����Ǐx��b`��,o���w�b �Lv��.c�:��Lɭ�$_�D���$�pL�S>Ij^�q���	�3���}����nf���P)3"�^S\�}�[Y)��\�ɆZoi���`����@�ԕxpT��tnm������+1�z����-0Q���=s���B"�>�a��
M�s���Dw}�c0`>�fvqw+�ZR�ͼ@��Q����>������\�4nr~�٧�(���*�D߅=�<Cs��|TAz	�j<<��tĻ��Y�<��_���Z��St��F��j����e�iI� �&�&}_�"Jƙ��1_\�Ѹ��pv#*]���A{��*21uaH�S���Z�f(�w�����$��2>ӿL]?�o���ar\{ʔ(�ۨ-�,�K�o�;ڋN������{LO8%x��Y+�yǀ�v�O[�T�4�v���U�J�4���(��o�5.th]����PGM�FG1J�N3���)T��IX(�z�A�t��.�ВqT��?#�1+q$����<S��8y EM�I��=���u�"z���4�4��1:��ގ�����+��$�fѓ}�G���b�M���M�$J�Ǻ���y����k+��bIr�[;8.ލ�F����@�= �Ò{�A ��3eJع��cV^�=�j$�;_vε�Z�Qg}ML�\�&����m�&t键��2���=;�T�����Y?�����|ބUC6m�D��j?"�)��"v]���A�va1d@K��Y��1��2�M��5�-�,5l�}��O��">�Y<ZJ�ro�'+�u�R[��t�n����La_�d|��j�Fw�w��Đ����f�9�\�%725��d������I�t�{E��nJ�fq�Hu�[�dI�I��"Y5r��	x�>��c�?0���m���A�3��T��"��G�YV�������)���۬��C��""�Պ��� gH�R��=���@�x��+eR}��yK��J���Ŵ0F�]>z�t�O/Aﵕ��Olyz-����+
)���0�}@����$Bm�>2A,=(]�-}S��6B�l������������&4��Lb�H����Ԃ�f��o�1�վG[Х��
.�Qv�VChֵ�MX��L��O��͙01�㠟�;���D� �%�����x��83�� ����#�N��9k$�KS8��؆T����a'I��ʼ�ֻ�qd6��L�D���M;��o��keϙ�jb#@���d����z�>��%Ng�Pn�2�T�O��ac���OR2g٧���t���h�Ǿw���*�Nz/('�.�!�u=�8��W1����y+�w-�9#���Zj?^� ��ù/o4'�����P�+���U���b����j�0��3���P{�TL��0-�_bꢢ|93nߑE�EU|x��?_u%�_����K&5�>�Y%L ����8���1�z$���aO�ͱ_\͚�h��}ASq��8���sVel��x�}
nS]ԻKT_MQ�4���a�.4��xa}�C� �g���ٯ.r�1���s�?b��EGD�#�:���!�DZSS�=�EѢ�NS�_�ȕY��?��K�OZ?$�YSX�0B+�3ʤV2�s4��LV¼��̪?AW'C`�E��� ���#���j!��MT%�@���w��ɤ7B����':�?��4G�܉J�{u�ɛ�_�E��bC����H��N�=��n�'Bo���%2�˟CԪK�Ǆ�e.���'5e�y�˪���^B�ϻu�����]C��J�����W�w�P����~�f
��z �w}?5��=N�'a���e�e�����̠KPA_��&}���ඐe����0�)ܵ����&�u댾J	�Fn�(���t�� ��&72qM#���.n��|��)	7�d�S��$[����:���u�y�De�!k̏��5�����p��`y�M@�_����'P��-γ*~q�����9�]H�ѹ~D �qA�.PN���[(;l�Sڶ�<P;��M�aM3��_�c8"L�q�Юi�F�m%.�N��0:�K���l��)GT89�y�$T���ʝI�"T%R������UB���A���Wgԝ�ȸ̞��빵n��T�����O��Q��6td�j�m}Fe�'KA��;J+5��#!��6�iȋImJ���=�?S�h��d"��2�z	rY�֚d}�ɕ��g�Zr��p��������!�_�$7}R���)x ]�hz�֨Y��_�,-��^� �5�=�GT��	)hr��O������DpH%��	�	7��j��E7����S�л	�9��J�$O�l������R�OU)�=돤�[{ :��ꯥ�
D�E��C$"�ߐϳ�f�y{�	�R������Ϙ����6���C�\�SXΰ��b,���{�������>-"R��I�|������~t���i��*`�'�j��}�P͗�1��^	����:��~�S����T�Ͱ�B�\"��ܴ��e�&�����2v���	��T��R;=�}�:��y�������z�7�z�zO�o�[���7���T�]�ug�p���aʶ��DF��2`-���}fɤƜ�>��\xW/o�OY�;r y쉹\��%�������M�}{\�T��_T�s�I�BG*�dW���ȑL4*R�Q�wJ�-�=��B����E�?����ٯÉ�5^H�{<817�"��,AV�,��؇�<�����m�sk�1�v�g�":������4�]��ǽe��Np��&ْ�Ƶ	i��2ER�"9}�8�=���KJ��O%�o�L���Ր�фG�$$��Y:�'%	_����-���t���n[���N���8�*�p3O�t�1.�|E9������{�?�q���J�Aй��'��לPeK��cѲД?Q�bi*�O`����<�Ac�D�\��^w�r�G�U��s�q�k(�g^�xĪ�v.����N#ؘ
��)���h.�d]_���5�b�M{'��L5�Ϡ ZrPύ��}�Dw����F�Wiښ:��ݑУCY"_��g����E&PH�B�/F�76'J<�t4�c^aKU�̘�q����!`Ȉ����_��#Gy��B�_���o���~�>�Ұ�t��4��0e|:�%����,
����'U)?�����8WLq��_c�e"f��yl�K[������۵�b�+�,��� t�?��nͰny��I�PYN���OE���b}�*4#� ��LH�T
���ɮ�Wˎ��R��d�!�/��*ک,^y,�|�K��*ȦL�@� ��2T��O5��� 
g$s@�W�Z�xߴ4N:2N�]��Sd���^2o��!�;d�,+4`qk�}�W�HR%e���\0#�^�ѥ�I�YF����DC3�u��R�`� >��_z�Δ�%� 7�=���0�u��>�c=��*�2�~p\̉|�O�ipճ���AU
a_��wݙ25��V8i�̐
�O�/f9Zȹ���|��HK��>�s��>�C����b<Ӵu��s�ϗ���Ba<"��T"�S������l��l���͎3�R��� �ʺB���g�q7w�뉨_���N�րcL�C~������*�0?Җ�׎�h�Ȩ�1e-Y����ulO<(RJa�P�nw>2�{f�A������ U���Cw�#�W��
)J��Cz2Eu��'h��ַ�ou|,?������q�ڏcYUhۏ?.*�u~��hP����OY>Y)̼S�V�a���@�^9�h�ɖ��)f�Á�\����o7Ss�;�?�E��=��9`�9P�k��r�I4�<�Fr��y������7��XlHc�-Kg?�Pd��;s"`>M����~����9� ��6��!�UH��G�*��I�b$u'r6>>R���SM��eg�dމ���$~�_��=���~��aC�rP� ��� �����z[h�-4�N:��v)�z(��!o�ͮ1���±�j{�$wd�@$���.�����HX6�ܛvnv��/��A����(_�/l���K�E��t�x�!��s�Tg�=X��X��Ǆ��qR������4�S���k����(�&fGh���)t/9&�(������f�$%��v�h]Eu�2��!������Ա(���wm@�wI�0,ud�BI�_�.m��x��x�����z�(�6��x��2�j��l�k��@�.�bE�T�Ii2��J<S��EC�r����|�w����7����f���m�!T�X�>��o���@���O]12�&r[Fn%����	vM�c2�r���;�������Z%�Ǩ��{	�����t�?�q(O�}��2����6�:�w5����2�Rk߭���bTK�|�qK�~�J�GA~��,�؍����V�Y�,~M�E���nz���`xn~�wg��~0��z�=��"�o�F৏����!L(n�8�N�E�unbH"ۻ�o�]B��9C>)�!�en�p��K��xd�,_����}x{h�&�e���kS�p�1J	
=����sZ�����,5��u��8�h����§�O�ïy��w�>n����{�[}�0�'gf��2e���BHs�C��:k��Z�|�ڕ���:��W~+'>'ˊTT;����7JDhf��v��rӏַ�֣�ܶ��n����B���q���k�翏�{��(^�%'w�_խ�S���� E�7(ԝ'���%�ԭ���?d?�G�j �� e,0������J0�y��:��س.|�b�����Ƈٞ7�DH������r_Cvɡr�
�}Q�;���8-��]��8���u�?�y��ܩS������f!j��f��yel���"8�5��Bv�P�|W`����?��c@E����a���=�>m� �ou�545y���!��+��bd�p<�3�f��\	�5ʲ6���"�#4��Mzz?��+���3+F]��a������g91���A�is^��'�Qף�.t�������3�[��\�u��\8�����`�+�v���R=��i�Cړ:zE�72;.lnz�m�� Jvqr㩣W�	����p�;����"���T���ry��RG��������_�*t������RI!��Ha���[�*(4Ǽ"CͿ߀�X�/��c@8�t9�}�^��!�)F\�ir����=�s��̰2������sS����g�<��� /?�,��z����%����<�&�:���|��-���q��Zu�,�
��"H�j��J���6�
O�U5Gh�
���H�a"qk��-�Dc��^T'�@w߸�5��
�]4;�9��}<��q��㍧�d#��P�W�O���j�#�x��@�h
��M�,z5vGyC�K)� v����Թ\�N͎���kc�ٌ���j��,�'~G���|�bF�1��4?d�2�*�C�q���� ^�W6G��Sq��-��kYUa����A�gV2hD_U&ކ�2�!��7��h�F��l"���^�����D��P��,L�G���\�{J�8�~P�s�*-�n���_��cf�=�`��0�#a��Q]n��ǥq�����#p�G�q<W�<\Ұ���t2w�kg�g�m��X
l1�h�r�y��d�bVDb�H{p�@2�J>���,L֝D
�Eן	 phь���;
�R��*9R���S(�������`;Y��N�Tc�"X�Ȉ	K+|�Ck�+#O=��Z����? ��>��~Z�	*m��T쪰���K�c��� f��MZ��k�(�x�!?vz?�A� ��/�U�̮��R���`>�r�c?�d�������h?X$��rR����h�qR,�Lv�=�D��Į�r����5����&oj�b�~�Rd-߯1�MM9�7�\� /��KdDs��� �n4�.��'�7�~��b��f��4��'���C�ipKrZ\G�ʥ5�s��^K1�)_,�/S���L���
��6����2���X����pQ�Љ��?�x�h?h��4��9����dS�b��(�ʱ\�z�-2bБ�?�n�i�J��&�V�<~W����AGVϮx��#���*��bbL��%s������j�e>_{M���k-UQY�.-MN��Z��.�,ܴ�z�զtSxg�s"�=:sD2�NS��KP'b�1�ͯ��[d�ftJB���s"ӷEt�JB���蔤�L����~���*++g��a�pm�G��/8g6��St����5�ax6Ht�������DwOOXe%%%���6T[{|2���������r���>M,��O��񢢢�b23)���!�@�X�y���}Nq`N�XFW�w�n�f��$�[���)��ŧW�r+����%h�S��ӢSl�.Z:�g��gg9^s�CCAyyy\���)�*��������;������?�o�X��.LA#���n�������zzz��}u8�K�HII���������~�����z����υ�����"�g�\�Z�i3OO�t�Z��+� ���:䙕����jj��Y�U�B7d�	��	�=n�jU8�\""�.���WW��}�6�1��37L�ۓz�[⣡��WX�>66���2�ȥ�
$�{Ⱦm����N��:i�����r7��'&G�V#�I������N�hm`�X��d@<d6J�3e�Ȝ�m��}O<О�/1�,U!m���ї��D��#�ёm��چ����c����ؑ_	>*,,�v�g7���ѫ����sSy�#��c�!�h�Zd$ń}���GѺ��#.�.:\�������N�3�������(>���\���{9���>��е7_I%�����q	A�^TZ+���EO����wvv�]�Q�(D@�Vk��5�JI���>���ƕ��Mٶp���1cŏ��\����\\~�����4=X��\Z���Q�.M�/�!-�Xч=�o[��7���G&�'r�	���xLb����`}�5)����	��:]hǑ�:9����ij�c~rr�Sa���U��!�b�CjBJ���Ϊ��Ӷt�P%o�ͷgH�q����(YY�WVL/Wlll�����F�"`3c��u��2�6cQ��oʐ ��̊��'A���՗'*\t7Г�R\��Іffb%ޜ���6�o-u�4�M+��+�)G���P�t,}Z�q/��"B�gg��n�&�ܘ;����,--u*�����k_�D�������I{�#���$���f�=�ۓ�n"`�y+[cj:����4t��v 
�Ë�:��?q�k�슣|���ve�cM~s3��x�J�˨�x�[R��uR���7�f�G��ʼ����n0
F�@����]��m`ᡍ��I�����sڪm@��`@�ì�)n���.�b�f�<��E�����ښ�������l�����?���vź�(��\k�^�x��C���<fbbڿ��3�M� %#ãd� uhzsy�����=�))�O1)Kz�>�1��S��&��ɑ�]�Ox��X|�0:��V�b]�j������􌌃�)���<Y�Vb��(�����Fh�FXE��b�/�S�-�����L��?�&������P����Tf�{�r�]-g�뛐��;����`�'$?j�e�wj�����k�>;#>.�w��~�%��/q�>)�����.l��k�L1n��4��b=?~��>>"��o�Zf�]wZ			�X�2�9ɒ�Oq����W�Z"{�Z(�x��#X~��Nc�b��M�,r</J�1N��h�]�x��o�()A�I�:�O#�0���a�"""�̔xh�&�.�Ƌ�_f��46����ፍ�C.,hep1w��5r
�N͑gs�����^7�Vv4��p�Z0�u$)�* ��5�� �<|3XSJ���c��h�ED_�N:l��/蕏�,���|��MÑ���r�hYvGHd0����=�|�.#������liH���)B�����w>r��#X`[$ռp�U�u���zD����w�ڈF���M����d� %�8�ɘ%�����"א;Vg�'���F���[
u��-`�ϖxS������$2N�e.:g˵��׌�s�lI�gy�wM@q4^�6xߜ��..ו�L��(n�o�h^�����}��ݔ����`+f_b����,s�Y�d\m=)Ҡ|~Bf�;�*�F޷o���}�(�c���|C��?�X��^{�YT���!�6Y�D}�.����ؚo};�͖ ��G&z�ٲ�&<U�j��y]"���I�b�k��S򾦘�O�A�_+J:�)C�c@c��J
�jsMJI�J�󥇅����g����f`ae���'���&ys��a/�$*�g���S�)gw�Q�j�R�e1d��М8�������]D��I���U�&�^���Vyqwd�
q���T��>����ĨAɍU��'/�cq%ʤ$Z:����Uo�Ǌ��=�5�Vca��ss�کq3�4[Ȇ���ƣ_b�)�u�4y����I�5tx�:�Q����`*OHd07� ��l�c�!�����il�e��{�0�Ѽx[5?|q�<�B999v��ޓ;z�߿��#�J������]�ჭ�_�kZn^�$vJ^�ˊߞ/����oo|l���FT�bG>�F��TBS,���f��z"Y6bX�֏0�Պ�|-�qQy���8��x�;,�r0�����af�(Jzq�26���չ݆��׾��鹸���@�H"��"�-/ǫ�դ=,�[�����'������b1z�Bt�����ȟ��ݰ[��,`	岿���B�Z��W��izԤ�柿�Ȫܐ�����_�}i⾞ON؂l?�O�����48�C��^dDA�Ǐ	:H�+��!��W�Ƒұv��S����v+��8��C��� R$����-ɴ�����Dщb��Ĳ,��Ƕ�<
R�k30��)�qGZ����k�K��i�e���B>z3`ӳ��ã��`���{�T�=��ƍ�©$��^-(�{��ޟ8����9�����xSRxs0�^x�n
�2()5ui�aO�ѱd�
�`��N�A4�"�)�|�UqQ�唩� 5,����K��'���0�J�:^��N-L��IA�[���e..�pYwe: �����@���}Pf�k���¢�/^�&���*0F���a	�����$�k��￥���{�NH��a@��d��$��n͈*NX����<��%}E٩��-���3$Щ�c��ނ����ϔ�Q IDW���/yOO�����O�x�<T.	�[s����t^��:|�JXc?��0Q��=�[g��%��������iD������wZ�SzD��0��9�R鞻>�oT�V*Sk��5�9��`������Ƅ�dj2���m%S���㕕��u���/K��Oƴ�Ԓ"�ݱ�]�}y�<��i��<����H��]/=���"��i7q�x���.�<},�k���6�{̇N&�7�n,�?��T�%�D�d�^�Ȓx>J�
'��#���l�Ia~/k^����N��A[�Ġ��f$���ݻ�\@���)a���{)�.+1qp��[.���n��{�H(��s{c��k+qVu�!���v��ad���}�[��ax�2����Yb.�Ad�^UDp	������t�urIFE���w-lQ�z��Do&�c�p����+O����x��-NU;�~��p^�������<N�9�� �1Ty����5̭4����%v0�R5��s�(�0_Ij*�s�LawB%����s wb����Q�G���`a����"�"�^Ԫb�L���GD臧�u�0}~m�]�?{�-�l<.�+���k{Cqی"/�bUM��@����L ~J�<�&oV���Du���9S��~GFHV��=w���K/��p��~�ܦ�Y�{��c��		�{>�����(�G��x�˒�����+*�]<<�ٚV�2ȚC��o!���u5n�/��aOw�K+�V#��IJ@N�$����s�伬s��j�8��B��J�@ϫ��Xd:�Ի��SI�ِ5w��ƍ�0�H$1e��g�[-�w�\w����nP�_�÷�y�|ďeI��C��K����k$`:��Z��g�+�S����}�����1�'�?�����'����ߝ�h��Mʟq�e9k��ph�ժ$��b�H��G̫A�h�����%oH�i�ɡ�IZBBaV�Q���P�)CAy�$N��=3��1�6������o:� 0�(2��.n|��ܝi�S�#����r�;T�J�U�H@��#�� ��{����R	tsL|��웽�1;"8�Y�3�m�Ӡ���p2�.�GBMcQ~�F�Ӣ��Fȧ�.�8�$���c�SC~w�۶d"�5>�$�@�D����U��5��Aԑ:?QG�'�Cԥ3~ "`�z�5��a*[E߾2f:�s�o���P.*�>������k�{�gb���R���@
��4ph��G�a�KN!��a&�����B�k�#
�e�,]��s�k �[n�~���K�#nǌ�B�W&>z�͗�B��5��	4���fPB�N���(�E~�:�\[��:�J��d#�.Q(o7HGί��OرC,}�W�y��4�(�%SS���A6�3���jY1�4QSǂ����O��IDݔ��ǄrA?-�'$����"Wή��n�=6��Y��񕔔޽��)}eg��fJ�a�å�i9�y�\"���Ͼ�]y�U��MO^a!��2���vvv���L@�bo��_d|��r��5��l�E�Ѵ�N�G�)�밮w_��{���v�^L�:�� ~�f�k}{���R���UM_?�#�����(1��j�
Ը�����a�KU�P�������?�_~D��j����b���bqY.|
~�a%.[��K#���q}C�A��5J��
ׅ��6"np��jjVZ���̬\�����]����O���_�L׌E��d��2�QxP�APl}���6�J��x^E�r
PNNN>�L��8
9>B��S4.��!�ۻ�������W��?����8�r+���!@U5�2���`��I΅#�w99���8]���+`���jFUq����I(��}��c���~8yG0�蔛�X<KillL���A�~05wK|6�E=�Xo�������ڻ۫�%���?6Ǌ������u�?m\��]PwW��6���ݏ���,1/��bWPaa(�zU�ZE%k=�������7[�K�W�o{W�A���٘�!�\�;ݓtO����baQ������@�K�b��ao��W�J�X ��Bņ��Z�ď�_4*��L�[������;��Kg��M�ݜ��hO윖�"���}?���!W��������h�t�OU�V 3��@e��\���׭e���"b�v�&`�h�/<?&¦��z�Y_w��P��Q�Gm���i��uViS%��9��A��w^0c�u��w$�ܯ_UܓJ5���K�PVVV*�w����|�6�A	dt`�U{[(�\��M�:�}�1�}}�EP�ʀ�A��c����ظ��w�'���?�R�ot������v|�?"1Ɣ�{�˧��a:ўT��ڍ���3T�)��=~���	����&Cw�K��?�н`Ѥdd��8!���G�u�������f� E������*f��ꔖ���Ќ�{�2�M�q�\��'�!N�K~~���Ґ3�����V� �������)�9�,<wG �߇����)��ȩ����M��kj�=��^xO:����;�}6Ӄ�"��\�=& �k�k.�dk�kj`��@^^�����CI	�mY�n�!��Ń�Ⰷ�9?�֒
M;#N�*��p��w�d$���_��y�	|3X�H��ABa�yC˕|�"S�^�Ɉ�ϊ�mHr�R 6�n�o/r�D�ncq��C������6z�@EEf�Ġ�SeG�[�U�6�����X&갠 ��
?rB�W�U�eS��������h���T��%���p�έ�NQ�6�b��t���		Nkn �`.��������Id��{�sx��}�^w���V(��a7���/,?S!�T�R��]�u/nf�j�c �M�no`�"����l��t�a=�ߍ��L�fCU]K�	`�B�+|��***Z���_W( �(��Hr�v���ذ#hps�[�e%ލ���?}���Đd�M������*/�}���IC�Њ�K;9j�����J�oc>؞mz��t��Nz�%d0�OԹ}Z']���W'	"n�q���{�� W�,2y	 �h�?�I�OO��\R:�Z���[��>�3 2n3}�_x�
 ]Nr��?|�C#&��������v�����|� ���Mo�,jx����͙�ϯ�����������W��/��;���2Љ���^��C�S���Pi�g�kPTK�Ѡ;�oQ�圿9��mz#�E�*��jaa!$�%@�l_�H2ٸ�Tݑ�#�P�x�������c��ZVV����������}�U���<U2��b�v=��{L��f
4�*�|--�����W\#�\�S�8f�����W;��ɆC�h�9�~(Ѱ��&��� ��#���DD[���ō�����AC��owɓ��=r�h��&�h���?o���h��T���������|�����������Ĵݓ���'�g
q�WG�=a��?j`��u�:)$0�d� �1����
|j}ݦ���}j�
�|�bbc#�2�æ�Z(������'O��Q�������EǽK�_x���Ֆ5gJ:Q�B�$��c��j��,�i�900��2����$�M
��(
��n�R\�����7ܣ��Q`/�Yg�^<�e�Г��� �"�9Ի��$�@ }��˷�_�c�G�A��],�g���f#��d�D�β#����`/��ne٧Y��W�?�c�������@����_%�@����3n��Q�ܿ�S��~�nV>�k�I/�JgU�H^-֬��#���p ��ۄ�i�wMlN�.yǚ%*83�b��drhr��?�7@%7��c9��j�Hd�0YȦ �#|
Ђ����?�>�lOV*؄56�����i���
�W�~�ͺJbX����K߱~�IC[�����\����<R����{̷�ߩ��̈́��g�1OU4--�\̤J/��G�"UWe{�ۇ�������P�B�U�j�}��L�����Ibʷ�����[��>�BN�7�)�r888�~9	f�l}�)����"Jϭٴ߆!��o�1V��?�(��,�l�PS���X7�~�Ee��{f�9��0��w<^�`��Ȭ�*&�d85�|UZN���<9;3�����:q���3��q4�T_/��+�x�PP�Qb���_M��{�g�ֲYX���%��5��W-0��l����Аb��W@b�SM�μ�kWR�sY��0�ʜU9����0�rҰL.�thVKu51`cbO�w�!��ޞִD�����5�s_I�5�4��۳��v��k��f��Ɠ���r�pP}��3�H��V�ɸqNu�&X����������Q��ƍ2���SS�ZU%+311�yli� ��ٚQI t"�PN���v�*t� �����`~�%����W��o�i�J�~���������rb�~{9ނ~%��^h���1�;�.=b��$v݅����M����.��V�
�D��։���S�~wڞ���u�P܎G����P���J�2�p�����T�JU�t_U��$!c��a���_���C�n�`�s7��Ľ�9bC ���0S��>(+��D�l7�]�L�o��FE|.��Q�z�{$�����S�Li��8,7WX��'��=�aR�� �`P��))�����(���B����e~I�8����:�;�jAanjJ�|ZU��������Qll,��c���_Re��?�K a�67��&���b1-,�Z@P�0���i�JUa!�(��8�.B������ma���uR�����������uީ�L	X�h{
Q��E ,�}����q��������ӺRN��&�C;B� �UPfJ������[�9^7�`~r�����fd�&�(*��+ݯe^ԫ�!H����6��Y��wvv`���8���Y��z�\�#���ϗh�N��O���5��#n�\N�1��yz��i���29S��0��Ĩ��d��<3i���������au�4>"-��DF����2�j�a倫��:��'7�o��V��kG^ �T&����Ȁ�_>�����(
A��A�yf�H����O	�����[4v��r���ν�H��MU򄫉���J����	\��IZikk���5�����G���NO	I��Z3�g��G|-Ӎ��w1�)�{N����kklJQ�|K���֬ ���!a��ap5r0?wX7׊�z��Z�H��7r^4���)7�Z]��r�����~xf�P�m����[���ȧ��$�V�#��I:��_g���D"�j�<wz��H��[��w6�
�*p�d�a�@!�[�J�?���40_O!,X�j��a�,//N�W2���~�ǣvU�do�s� �V]�^��V���r��`ɢ�R;�?��	u�|���OO���4nj��/�>����_��W˹^f���@X6�[߾�zH~�]�Ǒj�_����=o��ħia
�x��N*ILTԵ�H��@/�Dr�s}0�!���,`�����g�#ڭ��S����&_-�t/_��ת'���e]bK1|�x�4�^���̂@ r�. ϜuˉaFlx-�DE�4�mG
��#��y����,��3e]���}r$��e]�D�O�A�������y(Si���"[ŕ�"OgffD��Q�v���������{:-�tT�v*�$�(���SB�$d��2�2bd�R�SQ�,CIʾOR�u���$����}��t���x~z>?��k{/���u]ל�h�l7m�S��9�}~�q>3m|�f�Bi`:P-u@e-�^r�����*���A�¿�'�3���(b����r0*M���>��TzO�F�aJ��l�z\C��y�I	�7�H$�ۙLbֶy�18���Ly����F�ar��ˍ� �}�9q�:^�{����O��?��jr���.��<o���;ց�j�hw�C��`��q����ܹ|�r�X�w:�����K�����J�K������w�ؕml���NR�z�&S�j\jKN�B��it|��闧#�E������}�8���������^@v���I�ߡ����~��c�`T��|�>ˤT����!_��e�U}�J�����666Zc_�x�tn�)1�%�"nyqV~J&��K�[�G|$Q��fi��������瞄���!�p0gF��p��G���<�ª1�B?V$����x����/�;�����r�����m�G��=�{_�v�~s���'p������+_ˢg6�VC������S�X*�'s�υ�E�D'��z gBAAy�Q���e���'�UFb\�՜�p �m���wI�������͹�!���74lݫk�bA-&��j\��j�f>R!+�[����:Q�1�s߂����_p�RGI��+��}��
n=�'��y�Lz}=-A��"s�w~���A�l��ڴ��	y�xG㣖��H�vl���柿w�9�-�6�q��#	��풢#oLs�TFυCP�z�`��M4�y�����-I�b�Hj̼k�~-�
c�X:���y�+��Xw�rVQsrp�����A��]�n�qϢ��d.3ӳ�;�Hz���y�2DO�z��]��W
���Z�v��lg%�/��bMRsRvB�_�Ȯ�:����!L�,���������~y������aջ�P4��W����f��Q6������C���5H��NI����	�#�\�n����LLK��+A��j?�u����θҖ�BQ��QR��REfG�m�8_����\&',��Y_/!--�\��6 ��l'���7�ͅùˤx�g��D\�	����0ACkk�HGN��U�z�f̡�J>)�5�_�k�Ioh��؄;���\�|�d�*255U���Z�;KƎ�F0e�o��F>��dv4�����Z8|�s!�M���O��B5ك����%cgZL�ѫQ%E�t*)����Z�>����!L��˝0K�K�O	Q o#t�x?O�+$�b�/3v�p��`+���$�Tԛ�(uujM��'��]k܅ڏ0��y�����_&[���-��%�3��m�"cJq�D��Ϟ ?�suX~��g�DZ��w,y�d6�`�*���oa�9c�G�:_�y����o}n���"�}���V�Á�Q��0|QQ��4��>�y�����P#��=h��ڦ,+U��2'G^;�P%䵹Ր/oE���$�#�5�B��$s�8��X�>.������}�FS�ڤ���uסSP�JMc��\�̕b\Y��	"���'�QDQr�iyc%���ݪzߙ����nD?�g:��C1��B�k���w��-.,8C�#�f�ݑy�tR��|�S���o����ɾ���M����[���p�1���� U uE��,3���W0`6,J۞����GP+�ƭ.�3<��{�]��l�p�n/�"���n��Z��J?��ޘz���i==j�~GkK����zu�U�M��]����ҭ�'dgF�{��z���&�"�ɡX$6��ĭg����.��GcFGG-W2H�,�;z�niEQ$m�Xx�� �|�y��Ҝl$��///�/��HWH��ѰOe,�q����
��J��5O��_�9WK�(��l�q:�׭Υ��+��if������ԫZ�{m�F2�3X_O�Hb��'���G�:t]p,S&F��\��/+�� Aܯ
ۆAK�S�]ھ�,p���.YSw���~V2�y -½����*j�:��D>Hy��ʴ�j��0����8�ɣ��G.tֈ�ųE��_>Y�}�1�o�Qc/��Ʉim�R�DQ��C��U���ZC-�Lʾ"���%`cg_�-{a�b��4@[,3��\O�.<d�.9�:�Wo�*�y��o�Jߎ8#-�M�ЬSf� ��Cy�x��@��M�}||�+\�ꔗ�K=������i�;�*��؝㡼<Ք7�ݑnߜD�ѯ���y��Utл���Y �ǀ�y�rN��.g �ea m�4o���a�vv�Hf���l�7�)���pz��b'�/�}��%��)�7�w�SY(���ﷺ���k�/,�3�UQQ�U���|��Y��qE=���[�Ͻo}mBrr2�3��7!�5�s{��~�*��<��v�% �"�����g�����$x��vc��p���hfW���v�?�5Oe�o���H"������H�e����<~��`V8��u���r�7_�����s%q8�D �,�2۸��ҳ��\����J&[!l�߈�ظ-p\�}+���:���.���y��͵��kN���!�������㽗���Ͽw~�������)`�o^�_��u&��|x F+m�����~E�>�jA{m��v�˱S�v+��������荏���{=�U�16�z!���+IK�^F���>�l��ƫ�	x���憙�z�?�T`��KΝ����nd��&æ� w�� ���L�{)�qj�D������w����e��Bi|ak>M��/4?�Ij!���FSbb|)Y�<P�%SmQE;��s�5���jR�E"t�y.�b�:���L���&���::L	���G�C,٧E��A�Eɓ́�#y�kJ��}c�o` �X��`��T��l��R��<���TTT"U}<��˲�[��g�9#��?8X���7Si��,L�Qk[[$���sLj|�Qt����|k�C,qTE �������B�_���j]��l����,��u�R,�6[f؝�<�(��N��ݝ��(�t�9gi�g�#�)鶍��6��ϰ�پi�U��_o�N-:ţڠ ���&�m;�S�>l ��g%�AJ��6���2ɬ`n����OnN�Xr��װ짫4�	�d���׏�u;�����n\�r��
�Te3��к���'}���Ɠ�,uĸ����O|��V0���XK:�/���g�����K�-P��$�ms�$��Rf1P$(�ס��ﻍ�c��	P��XT!��A����CE��,ĔJ���g�N��$K��yU��h+��~RAAGD�iN}�,tpd�*pagF��6:%��B�1�ZP�����p�d#O��p���������xc�V������E2q�:Ɂ[[��X��?�A*�9�ysSS�N!����'�E2>9Y�Z+_�i(�iJ�KLA��{2��'�nnu�|���=��a7�g����6 ^��Q�I�\7A��^���g��L��gx{�x�@�8���hZ�%ۚhy�b�aJ�Y4V��H��;6�}Tr+��C&t��9�eǫ�j)j!p�`4K�Z�d�eH����p��y/�l��!E3�*�����R޽_�������^�s({�oDXp��-�����fa�h�A?�Y�a�"����LPR��԰�5���]�³��̗�AJT�x�����?�������G�`��?��XdҒa���M�;#a�i������L>m�k(F��(����#�dq���OL,G�����pA�%)�������>a���@U���+`��`�N�u�-�װF��0i�N��c �M����=K�=`k,�x�.�&a��-��Mt��Օ�7��ʏ�Z����.����BQ7���G�^�ub�Y�/�������UGZ���M���h���w#*oSs FnwH�����:�[��t�j�*�DH�Sw���;�� 
����V��4�#N���Z��C�1s#V��vO��O0L�r�2�~�,�-����'첆8B��l�e�5����-�H���N�ӎ|��g�z��5b��".8�lT�,�&f��Ϛ�WZ���P��[�$����MѴ����yA٘/�������2�d,��j�ԥD�,����0��|������ճ|�]�N	V^79P�e�c��l�Qm����o��S��`�p*S�rf�d�MF�AJ�uV֘���:�W@0}��c��f�����_'2�$(�N 6ɒ|��0��0�f�d~kQ*�M���fn��#���Q��B+U�{�i���Y%*S)R�Ù�0������0�:KC1o���9z�_�����^��)0�����{�ؕ�_�j�a������v�1utS!5������?І#���e����V����w���xY���)$������Ħu��=%yut��Tτ�P�����s{�ML ��'�^ddd�ݢ̄���B&e�4
��Gy.��
?|����؇{ܯC�ԇ������'���]���q�.5%��GC`�B{�iE�`���J"��t/vϾDus�k����`����z5*`�����B�ʘ&�#4
��tni�N��'�������- he�|-	겋���W��y}w���&�#t����\r
�9�n�iΌjE����_�
�f�:;8(_fd��<�d�1Mܩ&5�{�W0ٝ�JK��d�����񣦠gy��2�����1O݊����ء`�q�6��ܘ��L������p��XՏ����Ϛ��ǖ�uU�?�ġPT?U��M-͇�xNW��v�S�ԁ;<h�2��{�;Z�7Y%�q����oW+d�9h�~*�T�"��K[�:��K�?@hN>��9�m�����_�c��@yo���{{08�"�dW���}Gth	6gD���y�t&k4E��Pl.*�p�N�V��,��M�3�g��1R�A[:W��_��T��c�F��[]D�0O�����le��DN��TR|�>���q��Q����#�<A�%�<���;�����F�d0����W�M���Pݛg��'���^��W�;^m������{����yX�﬛_�nڔw,�(�B����1H:թ�\�S���+],!v�cܺ=�~Q��}��H��Y.�B�����b�\8.�w*m������	*��v��mF��<��:�a��!J�v���c�e'�V�@��d�T�k���O��N/~)��P�{u�[l0he(H�&��ʰ|��#�7abM�m�p��t��T��h`W�3��	� B��;s�X
3O$əihht/��k�|��B#��f�s����~�\Vy8�O�U�|d���T[�#��y.�p��:G)cމJU/�@�����'p+�����f�L���H:�}�3?���}�Yb�SSS�e���[�j%6|E��Ef^;�)����M�.���ބ���W�����/�t{�����?��G�>b�k~R�n���7&��8�q��_��%�����bU��ĤOALV���L�Ī��^ �&%�Vut�5�y=<4TΈ@vFZ��v��
�&���}���G?^t"��7�X�(W���n�9�l!8殑Z��e�1n@a��Q7�҅�m�m�u��b0�[��ï��5W��|����w��E��o �QG� �S}}큣����E�C�?����Svao���1)��	TZ�a��Ξt���^縡��+++f�>�d���}0����ڲE�(�C^=��UE�w�_m�dM<Z���:����m�
��x�Q��}����7l�9~b���;%hH��[JC�2/T@g#�v�~#��U��c (��_P���HK��?z� E}��HY��V�h��h��-υu��D:��G�.T\�u���� vd_Ŏ�/��9�n��G�3��7�Ƿ�s�=K�H�g�R���܍�v�/��GZOY����%�XC��	�4Ƶ�Xqe��A�+��]Y���N�o�� E��($b��L[[�]w�R04B�ǣ�������y??����y�׭�	��%E�:q�*,�X�s�1�\[��C`�6��9���  �w?5�#4G� \���1�Ȗ�tW�>����n��.����LtRd]Vw���Ԕ�/>^ފ����Z��	/���̴��39p�m��1�9�5�C���:AAA�Z��4��ey�$E}=��E��@+����{L'[\ �_j`IV�T�^=:��*p����t<��V%"�q8�d�8 �j@2��#�'�����.C��x��7ΰ��/a-m�?D�P`������S"�ݣÜ�Q���ܺ��7Ywn��l:g u�\+����B�\�!�^G��i���hrm��^�����%Gy��M�>��]�JT��|�u����X](�N!!DѦ���*�v�4utDO�&���ԯ F��TT;<7?S�g���_��O��i�����Xxݳu@�2@�!�����4cr� �	�'Ť���bG��<���T��wc;֡�$�I=+#=�P� p���<ԹFG6C]S�����������;�YNߟ��E��X�	��O�i�� p7޴K���nIA�	��@�&�P�jf@��}�-x�ou1?�#%����ڪEl�Ⴖ@�2�������3��᝻\[�R+s�}�B�+|1���R_[�ϰ����z�#"��=�&]�Z��O��N/W���%��%�N�?ߏ�F���r��3vli��q�_P#��iddv�LBY
dٍ*H���n/怔�"v�U��XXa����t3F��j�����k催e�,B1��
�{���$�3��F��������5� ��p�B�<0�X��[xݞz�23P��F��(��dN��A�sA*�h�ϕ\���'k�D;�(�[L3H=�4ūv3?�PMG)��$>\?�ե�gv �h���!Q�����ᢩ��JR��]��j�4��0Dm����|�8�6:3H6�X�HwhM�)J�&[�,��9[�2>K`GIӒbA�6�+^<���n�˹��^ڟU���3�5�9Q� �+ԓ<�Y�q� �ډ/�Ǌf[LI��A��76���-\�"v���ߛ^�HP�Y��c���*�V��N�6cT��@qu��"�휄P<�l�r�R���S�Uz�,�'#9tt1)� 9�S�����jO:�Hqu���݂�&��c�t˛-��,A��9�n/=�����ȳ��-I���s�j�h�m����x�g@����8��JUCWF�Gѯ�*K�ٵ�>�нҖ��x�w畞bTG���&��+�p������N�m�۳�L�L&�-$B��d���T����+o�l;]����o��I�Ga��O��!.��D�ql�J���tk�� "$l�K��]��?F��1�N�2&��51��b1_e�E���M��.S�!)��g�p
VA
1߯��_Y�T�;b=�*����~�K�YJ	hƯ����1%a��Ʃ��0]�\q��ʫ���t�˛���Ŋ6������!�0��j��0�ɾ�1	�XAF$;���@��5��A?̇ ������R.z	�p�O��i��ŋ��-����_��DCNZw�"~�.R^�+�	:�-�k�1ӮiRx���!�[�ڲ����x�����b�_� ����B�3�?q�3��C0~�����íi~+Ett�;�ۍ��~�|	6��Z}��:!��~-,�;� �<9�6Ru$��v��o[�����hy"��S�"�x�
���������Τ��#0z��*Ќ�BP��;��| �龢B� �@�}��鷠�*����a�'����r���qhE�A+�ԩV.!��D�<P�~u�IO���5�D��VU*�l�C"�Х(�h�rA73u�!bD��H�K�.A�?�j����i��d�v.�*�@���_�$�G�������j�ʃ�`�R+ou�=�(�X��lR%�g�D�ٝ]��[�\q�Z�@> ��9�O{.,.�1�o��p_ɏ�ހO�L5�V���<<�����+����SScc~+cș�t���532�ܼ��C��P�ֆETR�w��&N�J�"�u���΃��I�2L���4E�cy�C�8.K�b�V���t@�`�Y�6�3#�y>�ٿ��|C�|��n�pQm��K[l|d\SOϘ�>�M��`$x�%�-�}���C666�5	�ۆ-�_�
))�n����bRJ<"I4>�'�mу���{A�N�q��n������Dc��Rt���g�:�#�qI�T/ё$���D�_L�iN8�����@ �����ݟ�����N������8�Z�ġ��]����wϱ6��d�ve��E_-����.Iui`m�_��^�vM/�a�mH>
Ir�_���A:�v�-��$e�R���C�3{+��	x�-l���AoL���^šv����p�S�#s֫P��y~�&�a�ګ(7;R�l��{�/�߅�+���M�8�0�ڪGO��k0&:��.P���#Ea�i�^�
�C�QI[(p�un��,�)���k�{��{@#��p8�gq�̀9$�:��I�Ep���� &��8�0�G���;L	x޽0���}A�ᦎk�(�w��� 3n�8���|�E�e��!k�7=�b����rH��'ӳ����2v�i#�j./�*+d�?r�^��=������S�]����{PJ��ss�k`�I��|��:}*c$:��X���?�
��w,[g&�������� }��+����߬���ld������aSRT��=K"n�s��6��C�,�}�<�aRp��ʄ��c��o������s�G9#����n���VG�+���|]��R���e��Y��IC01���8�� ?� �T��5�%�E5��������ԅd(�E�-۬�H.�D�Gh�[���...^��Y��n���=-��
#�E���2���W/^�=ne*�eu�	篤!2�2ڱ
X&4q�DQR��*�7'k'��WB�����/�;%���夥�;6yéZ�g���W|M�T����zD(�I�C~�T2'�E୥�UG��M<tzy�f�S+��;����s	ը�v� J	� T&h���^�y ��]��U�59ˇ��@]#J��P�XkA@=�.ŭ���UƎ��k�=�'��ŭn�W���n]�F�>&�&�܍�5��~d�\�gZ�͂���.n���)xX���&������fi��2�6���u&�,��l�N��vy��n�̌���x�&}q7�"��:���q}�݀p'�E��58Ej���+v����S�N�Q��`Q(܇(XNl��^Bdʥ��Md�?��4�._���uS�T���]��d�(�C*�4X�β<�5�����������^\@z�i�k���?��_����3h�=W�_����n
u��ZS4�mJ�3�Mϓ:�3��r7���;^I�9�0'�|�=���
V��������=/���a�%h$���0��R)t(�R�M�
�,sz�n�����;�~{�`�Q���̛��R�O�m��O�T3cVl�����[���Î�R��am��'K��|�MZ/�͊T��+�3���w^�:O�[�(��%s�^�n��{���(�Yb��pn�-�A�Í�����\�_�Y"�3by+�ؙ\�����]�� ��B��[�R*+?�� �W{���S�"�<�Y���oܖ}��P�v^ h���Y�,��y^3�>an����������.������#���=~��q��XW� }F�(u���,�u%�U���/5��+���X�L����gֺ2��pa��x����z���6d�ۻ�=�2X�����Љ2�f<���Jn�7H�/4�!֗�b�;-2�3)_����͓�(n���,|\˂�-�
���u�&�p�Ѥ���mzC�jx?�듰\��D�tօ�hOv8��|��l��4���(G]�����,|�3�e�}�D�@Wy�#M5<W�?ҩӹZ���ԧ���>��Y���;�m��}Q���	!��RP����jRO�O�˫��Xzj0���#�Bwߣ˰ 
�ȍ'�d�R�1��7�!���#�At�̥(fu����N�s�1�q�s�.��t��q��"U@��F�_֫.^a�$1H!��o��mr��uxt�.XT��<� 0=ҔHR�vU�F�B
�U�wR9����f@k`$1k7�+>���[�Qt7�<�<@�J�w2�JW~�������N���Y]$7ۣ�<�1�U�h󲩩I���2 �ۺ�]���"R��ݮ�m��/H�¯� �%޴�2����D���6!W�3�ۍ(/lM�=JD���ۀ�BB�Z�SDҴi�{��y:�=��9��
�"�&Pme�G�1�}V>�� ��'�-ۡ��j�
��h�GfI,��Y��u+�|�[9q���� %H�� m���n�b'����݅��0�2��mD=���е~�3#n�����i���=�뤈P��s�p�أ!1��Q�l��vRͩa6��d�+���B�S(�0��p}J�/Q�~6(�6���V,���t!��#'�����.��c+\,�>jF�~6/L��<|:�9�B���}1��h��V ��!4[,\�X�Ǉe�`�#�U�=�;�G�����j�^��b#�yGƯ�ۨM����G4]�F�7
bl���?)��Pj#���&��������[Ո�_lG��B�9����	����)'U�B�̃�"8����4yXo�EdՌ`%���Yn�MƊ��#X�M"��T_o�X$�\��O'4W���~:��d5����+E���!Kƌ{����/	<QӛdO�w�x��������G�LK���6B�R�g� �0C����XX;%{�`u k��$�jyB
5-���|G�Ŏ!�.�ɲ��/���??�Z4nU<O��ͬ����������1�v?m�(�`�N͙PN>Ǒ�?w2o_�f�� m��v��&!2o�x|Ү�g�qD@�*�h{}��91^� ����	�S���u������w>ڌǿq�֯u ��b񝓆�`�����3�nli���^�9������3"b��rFUK��j��#��X-.'�G����i�fm4Cn��eE���վ0�H3U�Y���沓����,r�*�4%iW8F��Y3'q�����
���(�ց�|6U�R^;@N���ڬFިU��x��O��,o6.�JV�@{%��^�/n\?�"2NB��F�ْ�NG���/k�^��(g����vz���q�~�����t��)�^�L�0��0�+�����m����O���������z����8V�3�6���"�ၯd�dY�L1D�N��<k�6����bR?V[�1'�s��Xc��hqzrP�'A��f���Z�6�]���+�^�vD�"��d����`��>|�6�I�����f�N�R�B���t&�Q$ڝ`�-[��hWd�H}8��<\���J���z��LY�ok��̗�y�	�^|,�>�.���WpJ�z�͒"���cZ��.���/9IU�F���p����|J	]cc��.-�K���}1،�_���Kբ]�R�������\z����/�|���_gt �
&z ��A01��.k��ϒ��{��6;h�/�3��h^y۬�5�y�s����}��u�݅k#i���RK۳�]��5	?hM���^Z�RjJ��4X*�����3�����!��t����͗��n� H�������5z��|{���E�>w��﬩��&�Jbl2�,)�b�� �b����>}	��2��f	mV1Q��T5�WD�4U�2c��'�Ӷs�a��3W�5(�V`�mY����+��!����9FS>�&�<�*:߅�oeufԼ����_�	�?���;C��<����Ή����?{m��ǭ/�:t�������v܎���I������m/R2�cV�f%I~�c'�,�����,��?=��P��G�>�L'g��"R\}˛F������
a�9G󰨇��1='��7�c!�Q���=d�^���f�z��؇BǃzU��}�_��kT��3Q��ᄯ��f���y\��ɟXD����B�=7=ؓ�ĲH����ԯ�4����<ND�H�lؿq=�W����N>Z:�~��C���bfk�O�5K��-��.j���Ekc����������-%�4�*uK|�q'�.�mp��5�I�h^hy��yUR.ӏl��Vx˛�v%;/��c�3pqx|<BMHy�g�w1���u�Y��3�m<.>>ި�� ��ΰ�H�#��[J�o���#���c��<��a��c8�aGkGGGdm�ɱާF9٪�U~��ܧ�m���ډ��gǜ���K	6Oܖn��������n��{�'�2�Nf��yB����o�PK   W��X8�w���  ��  /   images/805fb750-7b5b-4a1e-90f5-2022d18e6d35.pngt�eT]ݒ6�qww���=����7���N$xpw���!���s�����������%O�ڟ�eP	A ����*�A���#���'@��,��)F��A\R&�	ܥ��՜,ݽL\-@^^^,6�vnf&�,N�V'�� 9HNRL�;�軗7��@G��#WX���&$2RU=
�(�h�OLR���
	B�X�*�>�z�hP��2���H���;�G/��Ga�������0UD#�� �|y)_k%�E�	n!|�Q�xH��:o�'
�󊳡k���AV��Ehl�atܽ�V�}�-£�z��4*�����R��[C��sN,�4����t�P��P1�s��k�a��[��9Uӳ��$ceoZ���Hd��nD�N���z]`bX��;��n>��v���*/2��Ю+D�Ѕf2g��
ZU#��*�*�Ɏ�$�r\�gq+�R]�P��blz��r"�V�m�BO���N�J�Ӕ1>��Ptǟ��.�;���r84(#!*&S�����C�,�g�"��oá�l�mI�b��k�}�*[�:���rF�չ&�!O1ogX���@*�n��^i���KtW�U�,�p��d��v+�)tpʊ��мb�!�2�L��uh<�V?y�M P��<�	���?Sby�J������Hb��<խ:9�c��Qv|З�͉�c
�:���9�	�(���)HBOT�����p-��b��A�Aa���b��HȣqH�_�ۃ�#J��s�'��L�	B�r6���ul4{��x��i����=8�O�\QF	A�|�&�
>�9�Kv�mb�U��tbDev;ORq�`�o�Y����v�G�P��ˡ���h�3irq2��[�&�����l ��E�lP�骟Mߑ�J��2��E���b�RE��/��m�*�t�jz�Ƞ�*�M�'.a�+F0�6@��.g,S�P�xZ ^rߍ�!*���,�)e�q}	�z�"y�L�bTtE�Bs��$g.������u⾂)c���.ȉ@�F���t�>�b�XC��433�024rQ�I��ʑ��������H���L8�X�o\�8�qgt�w�t��|h7��*�� 	�O���bcP�����?y$S�>���Gb�gT2R��dܕ�u��|F�S`��Gz��)K�jY^��2��Fl������\���o\��8�\G�!�1&h�A�����m�"5��#��
�A��x���+n�<X~&Aڷ�cQ���V!'�졅��rx��}�Elv�4{↽) ����o+~i��K�#\�o�XF#��`�kL����0�TO-�;����"�Ck�������G�f����`b/ ��M��vgC�1|���Ou+�����ܕ�+nR�Q�1�.��7 f ��̫Č_��zE�E7�bc��v�ɑ�*�j	n�g�_&8s�S�J\Y`4`��J����g5%e����5�
D�6'9�eS!�G0���s��s�~�ԗd*@���%	� �[��J���0��)�nV���ݪ4UY$���G��6)���Tư�:�&�X?Ƌ�j����^�bs�7ߺ
J�M�i�S�ZV�:h�+zO�8�֕e�8DlF0�}G�SM.=4)r�1Mw�7��S2��Hb��)UG��>b#
��+0�B��6ϸ�������Y���Q�I��F�b�O��&�Y#
忶�&�A4Պ�@퉲��%�̇���5(b���(����7_�,�r��w[|�6�.$��W["3-��������'27DMbɥGg"yS�&�A(�3`qe�Qѩ�,?��ol
�Mb�KN�P�B��L�V���]Y �@�q"׬���p� �Lg�6gn�::$���/n�(��SʒĴ42��FE}VXD) QJ�|� �7�J&tQ��F>m�wzȥgg"��$�C�5	�:4iF��6/�$r��H{��3p�H�M���T���n^���ռ3 ��'C�h��GT�`�i��m�C
F7�;�V�~_f���BV�?�䪜B9����[�Ҝ������B�t���a܅�oV�ҷqi�t���a؅�%۬��/Z�-����:�B��/�֨�`q�{`9���@��"�k꿚��]�w�����C��0����$F��}�I����·�T��Qs�6M�C1��sX�n��V ��M��Bz�5���&�"\�/}Oto��#�ŋo�x4�3SHI��oWC=�/��@p�r�5�4�{f:�Yᖧ�d"�r4+���({I� | �B �!�{8��;�>��X�@;��Z,��l�qp�.����+����VR&���T�vL�Ц�ۅ���N�<��ٗOt^|g@������s�<�
�K�\�*���VT&�̿��,�F�ㆹ�-�P��4���:��Hy��e�=��f��Y���Vκ�f[j�!�Y<�&�}�R��u�r������V�v�Rݩ�����Ue�Yeu �d�R�{g`���y.�ddd��H��=�s����=q8���^�"l,��R���FJ�@?m��a\��-a*��T*ӛոe�:���:�
p�Z��A�f��T�]Hj�b���T@��1 �ah�i�d"�������3��h����_�|x���o��D�_�Ə��*>KR��뱖CJ�$2��v��fX�4�S}�Q:Q��:pEsR�#c\M�5�2k�̰�CK���������m|+'�dQ���^�(�r";E����;:���E�8j{�4Qsz $M�G�j�@�ä9�ˬ�Y	�׵�w��z�׾���>��h���;�Y'�(ݕ�Q�1gJ���,7f�O��g<C.��$d�� OǋG������Rl���f\m)ts�F��O���s��֥8=�҆�w6 ���]s�6���>�<|h�^��>�R�7.`(��a���gf\�����Rl"�V�D�J��Qh�1�<��֊̰Je��8��1�f��<�mUEH�'W�]er�X�A��hv���N��B9��vWC��i���N�12�X*�f�J���.�����ԩ+��N�cN+��KG#î�t���%��5T�����?�t�$CW�n	(��-�z�L�OѼ.��ƕ1�������(�Q^(}��v��I���(/�-c- 9�?y�]��ha?�R���+3����'�>ﰸ���d���z�a����^=�,�k� AP �W,��:O�7dcrP��8.^j�9>2lh�1�/	x����V
ퟛM�J�����.}񈌓�A"� �0Ɂ�^��U�3z���s������
�7���L������.CF���*�Ġ�Vc�儬vݔsZ��R$�2����`��3� g�)��� 敜�[�����^�3�<AL�J��r�ވG�G�>Ձ�ߴ���l)O�mJҷ,��v� >�z.Fe[$o�s<�F�,�xL��̾����}}��6�q	5����%��1��ŵ�4���=�HB��^%�m�������ԫ��~��ch5�՛�%��YCY펈��X���]�łM�&�"$�,��?�E��.����)��V���4R�\�nӱ�N���l��Nz�h77DȚ�����>9ѫ��߹���F��|�Q���ex!��z*�=
$��_� �y�tʹ�ǈ�Q�L	y�T�sNi�9��Ґ� �yM�7��)O;���)�̲�߽(&'�������W��;f�����=�`A�ivj�=KAͻ5����t���-P�G�:d�f`,��y��Wߞ�U l�x�;Eؗ��`c��(�q�ÕL������Cp5�7��q�E���4�e��F�R��P7�ݚ!U�h�Zz�c�����\���c��?v�cm|��������b^�_�zG��_���5泩�][5��q�J�.VVˣ��A��Q�~F���5��������+�,y/�N;�C1�XSLf/&�&�}��E���V��`��ow6wn��vj��ߚ̳ 8���[O���lԼ_F�%m�[y�U\��K/�u��FXAξ�S�^��xA��F��;��Ki�M�[U��۸#��j�$�mE=ul���Ҏjg�2hɶ�cA�%��eO���ǒg ��Ӂg�����U��մ�*�^U,�3g�{i��b�[����CvR3)��,��r{��i�S��'2�'�Q���R�>��j߻]��
���9((�=7�g�'�¾�V���BJ`^���#�J	-$Xy���	8S�wM��d�0��z�K��}�d+S��}xd�&��mH���@�0.�6�-ǭ��5�1G-,g@��s�boF��g��.����*D��+�A��P:�a�״f.��f���i0�!����J4�BM����JZ��)��?Ի� >f1ev���؜	R��؅l'=JD�6�lFnT��`�oщv#Y"#em�>���ə�*�
��UM_�_�2�pSC�Sx0��*68�]54_��� ��T�V����V���:�>���&L_�Ru��0�,�Ϩb����k�Բ�u�w-���X���Q���l�?T��S�bQ1#.�u�m���@�T����|�9��7v�ޣ2�P	���_X�/�R�j"�O��Q�����A�k�	)i�gR���]
�%?L�{��g���v�x����ZT�!5�%+��ɿ8�Z�~��"E�UW��$ ��+ʊ1�tw�X '�A�=�b�B�Uٌ���xl.a������|0	���	��G/S"kCax@��8�*�c���C|��	�z��7�7����� .�M����׽/w.�}�$���U�y)��>��US�PV�js��qe�dy��yo��<���L��F��E��|Yj<Z�b�z���0o*��O�Ƀ�4P;�v)�֒r��FTIw��y#�s2�6�N���"c��]ψy#ɟ���b���٢/"�l���۸����IS�0����a:?��B&)bl�M�<��pT?G=)Z���#����Ŷ��4ۍ�l;tXW~L�/7��볝�ϩ��t��_�"c; �������«�_~�_#�k��&+���>Be+�o�!mX�rX���x��hޔu)���2�B��H�ĭ�g�uë����j`��R�X+m��צ[�ւVǫ��:<�p���gtU_�(䋎��pP����}nMIj��?��L�A��n�?85�2�?�#��WQ1:��C&1�28j$�{tx�%&��\�8fvW�<�)$�S����:������?��S�h��#mx%�s���W��9�K�w�j���m�*�� J2R��vx!��!]���#敗�緵�Ƿ�����}W��o�!�#�x��/$�eX�-{H"�UܯAJh���<��hEq��;��OA~�]��0��ĢB'$9��j1��h}d��8���3���šg�:�c��W��[�A�$����}��]�����d��_?��"�o��O�y[�C�0�������Q���+�^ppMu`��7� hH��������������+����J�ץ!����M��'��H��S��?Kϐǻ���gI�1�kՋ���B�b�u�8�4R݈q����#HM75��Z���M7w��F�5���͌Q��^r��׫	�m�v�i���93�Ot���_��.��ٟ��.����8W��[�ǘ��(W�Df
��R�Ո�gL"C��v+�Iv���Ý�x"�{H;��l��9����R���`��ߩ�N��y|o^��ؓ�EҪ:�+�#��ɶ�
��*�K��Q;��8�1x��YU��B^¹���yR�a�BA��/o9��MqxW���>�@}:T	E��M��n�&��V:���g�_l�|0Q��m*�n�&���2���mSeR�&�cx�z����	���6�Tx�S��i��=���?������O
�bc��0�\8���L�"�ˋ�n3���t�O�,H�e�H@~W}͏��P��V�+�T`xr)�TOLb����T\���1 HWQ��ʃ}��ԫ�ŝx�1����y?|'x��.���٨�+�P���z1.�����>*L�,쯅�$~��"]O��N$���p��u����"NF5{�Q�m�O������MI����j�d>�u$9��|g� �h	�}����,-�\m���\ѦqV���M����/���7n'J)��Ts�w!�S�5��aE���\Yr��*�<�'O11�Pc&��ߜ�
K����Ǝ~��NB������Q�����@uf[߿�W.�`���Z�⤀�L$:����m��O���|o��{Ԣ�""8ȃi�M���á���wm������c����䚩��;�tr�e�Į��T�q���6I'� �4�u����2 W�rY rSin�����_9E0���4J���	v�'\5��N�ˠ�*�3(�� �Tߵq7F����B�'^-��3��������ej��RSv� ��>���o�M#1���|#.xmon��0=�3F��:�PE&��^BM~�������T7�&�fWr/9/�1�m������e�`YK� �.�k���0��]�+�#0a��V2�ZBh����#�cO��U���#!N�`¨�Tu������]Sܽ��K]Y��#�7�?N$��?����W�IT&Ҡ��63�j�yn)���$}�><熶u�ߚ���T��.���;7!U�
c90\��mx�.IM-�g��k1��w�v��7e�[��TL:�����!�+:��i3���8`�f��M&�VH 3�[�d��$}̯�"�, ��#w�ϔ�?�bcqo�)�QL�6�2��3���jԂ?�vk�i֦��ja�IM��qb������(�$P�N���Ŧ�J�w��M5�-p����?�Wd�C�o*����ȝ%��3�TjJ��f|5�m��,�T�w+X|x� W7���*�C����N.�8
T4��}�T��	����6�+yg����f�z��T�/���*F-zj��&sU��/��3I,/��)v!�|�ĺ�t�=�47�bj����k��4wv�H[9<�1�ރm/<�R`���T`S��c����b�3�����L��4�	5-��D��� �e�w+z=��	�N%!���N����j��%�r��O>N���8?�)��I,?3�d����K��j��J#�<4�b�h���L~��S
��\��v��
-/<=`4��i��7<l�*ڨ"R�,�r�UFU���n#Ü���k��;�D<��A�����j��} e\@��Ж�R�����Sh�lzU ��t�jv�ۓS&'�V���d.�	0��ߋ�o���}�H�c��ešA���i�U�����C?O'�ԑ�Lp������r+�P��5b3��g��zz���5~b���`���q���I9q�}
l��J0�L�r]E�1�c��᪓��?�=��o�OzU��s£�NG�v1\D"6E:���a�^X����D5hU��W��L��s�DV`�0�r��-p�g1�H{�@��]t���T�� 2U����5(gd@����K�*iL\}G�"����pQ�2l��+}&�Z���9lݠ���ʑD�|�Uҁ��[bed��Q��Y{ű<O �FU�:��	�?���c?��T��*�h�,I�@$7�'�eɪ�$�XL5H�����2	h�8��?n����o���Lf(�o��0�i�8�pK�^�����ȑ��sa$�B�;�?s�*A⃗�,����ݓV@څ[�(�!��wJ��|ğ����3���o�6Y�e��&���cp}��~�#����?ҵ�"�&�*��fETО}��tխ�Dq�Se!=��M2[ĉ�����k��]��y��64�Y뱱�p����������3��A��f&�\�$J�YOW_]��#��ʏ�t�)�s��3}�-��eHM�]�?�-��fkOn�M�J09���J�i9*���Y%�"��䵂ڙ�w��@wf�A|��x����j�H�rn�j[*�q�l���#jzS�B_��U���T,w��`�OM�ٻN��pC�C���	I:�*�,b���:Y� �C��<��PQV�=a��|'�<�B��.e�����a%�i��2w��]o���>�{�S��u�3�1�Nc���){��把g7�p���̑�	�B������Kc�����2�ʵ��v��[��'vz�#Ó���}8DÚ�k�z�1�ᰐ����Yko#nc��L���I���%�����h�v�B,5X���%���T:Ɗ���H�u�����p������!��r%H��c}�x`s�h|���ߓ��\*ɰ���Jl+��c�@
�|�z��f���-�&��]�i[L�!���`	���q�yrb��㘰�Q�C::����r���l*�!%geЧ5�f��O�=�;�mC�ެ����S_M�J2�����(�k�#�Ō���t�3�%��e�WG��
<�W��_U�s������c�k�.�)��'m���n`0��U���i`���/Nmp{?��g��no�t��\� Ǩ�F0����x�B8�O�B7;!&Nx3���1��
��>�U7�R�K�����R5��w��~>�%_��`�G���(z�m/-��pC@%��ij�H����$�E��OFH4Xj�J���A$���k~$�e�}&|3.�G��ʺ5?d_�{��z� �<����z$�\-�si)s�`v6_C�p���]^-8��h��yzv��{�[e��aq}���:�wvgW��m~�?l�do���ZN�]�ϝ/}�x�����ڵdM�m%�H:�7ܵq)h�MVk�>�{��t꽼�\"s.(%WLjU�j�֥VW�e@�K�9ޙ}��'�	f�|���-����͍���(�Z�s(�r�ӼA�D�����56v��9Ͻ�YMڈ�-@h��=�(K��$|!����]ܗ�ά����n&Ґ�`�I��~R��I3�ý�j�'^N��,��E���ƞ�I(����	"��� ??�����v8	-81�/�̎M�sj�,p�.���d���O��亜�D8f�����fM� O,�� �GAUϓ���4�2�0:���b�`�q��]O���]�Y��`� �E8�{��S��Yy5��l��e�)Q�I�։���3��+�b�{�����3��fx`lltY/�A���������zW�w~�Y=hn:��፛?�b~d<��:��S��u3U�m�U��G���������A��h�� +�~��*�F��4 ����J5'!������ta������yn�
e
�0��62�W?t�oQ.ѱV@Vn,?*+�c	�s��T)i	�����"P �{�-ݜ�c5e��F��{Z��mﻡ���
���ۀ L;L:O���}b���oa���{j�ߝ� ����dtB���eѼn7��pM�5�����{���Hd���l(��`�A��LBQMD�F|�iw���i��-�b]��͂��p��P�nY@���cT_�.Ywo�������jID�bh�y�Q((��}����h���}��� !Gۈ@�ȁV���C�p�0πɽմ��j��{�[�Ht�m4oJ lŘ�Ǽ�T�?�*^[de%y>ɐdS;&�'M�����t �W/ט~R�~�k��%�؛̓BDT�l{U�<�[��%�����i_ߩl
��B��E����zi8=kY�v��$�K���|ۙ#2���dɳ��i����@���;��� [L3À
��&��ۆt��5%�e����c�~ N<T�9y�Vo=+X��Ei���g#���\�d�9��Čp3�ݦp}e�3��>}Zy�N��z2f�m�c�~��aF�>KȌ��;�Κ�̘ؼ����c`H�ҙ8d��	������e����x�#�l�C`6�Ҟ���mWge���Z�CPu>ts���R�%��Ȧc��]�W��==��k��0X[=׮ߓ��N�|��+�^b ���o�Z_G)�3W��j�92�l{(詭��y:����n<���&{M��acpxHBE� �P*�&�����gO����q�%9D�Σ��
^:�1���,e?���LwCM][��iwD�v1<r53�$u>��BU�ҿ��_'�$\�R5�9�v5�7;}w;�m {���[���G{��nD��-���l�^6�:nj��ã��7�=��[�݈��ib�IERCٱJO�&�۩�.�4�-H&?��7RK�-����w�Ԓ�c�����(B��̯"��
�������Aۙ�0��먝���gdЊo�	�˪��U����z�·����c� �_\�k���c�-�2VpC��e
zo0�����1Ds����s^��Og:��f�h/�[��xU6���#���޼��ɞD�-'/H�\��a�l���}I� �G&�j�t�sK��g�bW��\#�=�� ei�΍��4���� Ʋ����VI(����u�f.	����I�����k}���ʅ��-�v�:��I�Ѯ����<����x�=�鰘#�����l���6�js���T�i�N"��W{��j�h��+�ox��̻ C���)ѓs�E�pzx�͝]��q��J��͙��{j�a���j��+��l"��΄.��+�[��9��s�*����P���]��z�s���fu�t��'�ZY�5��/4m>��$�.ӎ��`���{'�ǋY~V�R؛�(��O&}��g����N���ڐ/6�v=f��(9Tl�rXQ��� }B>�9�6b�sd@%��� B���y2W=�.^�^Þb&�^ԫ���Y��ؗ"�h�ܪf7�I����d��l֕��t���?�3��8S�����Y�󭆊��x�^pNJ����1��Yǂ���1�:s~�������@�����h�a�b��%�zh�a2��hOzfl���G�e��ӟ�e&�58��Z� R%v����-���$�O�_T��s�M�e�>�{���{��Q�7��h�9 �>..*✕=�[j&d�7bz\x��P��r$�Y������Ck�7ڌ��>uK��d��|�6�ǯ���������q��L����9Z����q�j[��6�.BZ6�_��\�� 0�콳6�������;�|�J������}y̞ޜ���ޟ����t
����Vj��'a�׈�BW����=�@|k9�4�W�G�,q��n��~ӺM@���~}v�EY�΁@�U����B��ŭ�AY��―��=�Ps}��V�m�E�3�����H@�����S~~˄�4��|u�խ��-�����Q7�L�fTE\�|9������� �*˻N�@�)��
�|�+˔��x���P�M���\��������6Na;���ĵ@$b���d��q�7n}��1�^���cBW�y�=�_�^絶����*���q������� ��ǣ�]x�� �҉��Z�>kN����2V��%z��d�t�󅹌���Y�ـd��<؍//�Z���A���v;�>-fUy���yz+��ܾo��sK3*���/�&Z<6�S4:�s�U�V;�����<�J(&MF�'_��n�&׋�ʭ@��?i6�������nk 2�֤�b3�>��
\P�\�=~������>�DG;X���O{E>_ �
�UV��@j�m�A�����p7-�������GY�q��^
���?�n/�\Q��Y���ڒ���|i�"C����/� k�C�6" 
���9�N򕡕	�8��IZ�x�iO��G��0gD���
@ț��޷@����^h����B�o���v����S&����!h�]�" �4i ,[ϐ�����{Y�qc�&[BA�2X��8�x{�!<H�'�zά�G
 4�;�r����� 5ҷϘ�4��j<y$�ueB�w��P�ԍ�p!&���ߓ�<Jb��^��R�ޏ'l��P��h�-'-�)�8]M �L4���ͬ
��?u�b+��q���o�̑-nAy�K#5S�a,�ˁD���鱃7Y��[�=��Lޯ��ָ��h���L����ۑ&q�}�[݄ɞ�Qvv<T��n^��&JF|�r����H�����Wr�;�h|��"}EH"r&�0H4�L~\����
��.�E,��v�_<��9�B�Q�8����J_~%�P�n�h��l��e�����gN�,ը�
�����.��w�����5&s~��P�P1{�7^�D�v�����P)����C$�������:R�6z5$<��!�~$�����h���[S��y���Upm�JI\��k�6�f��A�Ɵ���vF<�?��;�q7L�]�M�1��b�R������ŝk��V3���WR/旘��Ɍ`�jQ��J:�t�$A��[�8�=��<����Dc�z4:���O�P���t�/�>�.�ߜJ�ޕ�:��1�d
�i�a�,�����3�7�8jH{�,��.��=�v�GY�-{�ޏ���~n��5��ΠMN �4��z1=o���m�ZG�.�l�An�[������`�!v��� t�0P޶y������{|;n�
v�E~#�����-���4��[�?IO\�X��t��S�����\p��oHa�t5�b-Էd�u��U�:"�4�>�t0'�Glǭp����<���r-�چ�p4}�<a!��a�|yFu|��K��N��z�  ��n����>:Z�ĥ���b�M9����BL�\�������#�~ �i]���]8�ݏ�:r{��y�eN`f3{#ާ+���k!����U&�Lа}Z·:�5?Q0HqÞ#ޗ�o!�]FU��8�5��w�TqKq_}�	c	I�|R�D��&��_�l৕/���Om��w;d��0�wfKb�����y�(�(u��\��u���Fa�������L�A�\�_��jP�bPihX����k�!��I�y�eA�9�f[j�3%�_����M�T?u�>��ru���c}/:Bz��Q��υ3��=�4�d�g��0&��?�>m���FȌ2[b���6��6`���(����^8��#���l������۬��&__d�s��_��ӎ�٘*���oI��8M��,����i$�5#�#�� �c��,��|A����2Oӟ�&�'�6��,s���z�����/;�G���.�Y-d�}VHYݍ�Pg�Id+q�Q
�}���3��J2��F:弜�z;�yVU��������.g>�u���@�;r���L����,�ɣ�DԏM�Z;��F��J�IXb���cS��ɍ7�*�RX������+�X��Y�_��a����������|xg��q�7�u�c�~C�eY����C
�]@҄7��p�5�4���]}��lɑ��
yv�\GG?��fz~��*�Ts��x�
���u�]�k�W��Fч�	�Q�������W��׷h+��M�hftK�3<���S����7��|!��~�y����bIc� �v�w��cb�����S�J������Q�������X�Сň��XI��퇇$�߼H���~� P(u��q�������T�L����9�dm�ë|fUr:Q�QX+d�^d$���B����QX)�q�G�+rrr�J��x��u/�}[��!iD���[���KQmt"�Xͣ|��5��]���~�^nc�u��l��c0J�o<�C�����E�k~	�o0嚱{E�>�L�Dp*:j0��_LE>�Fq�o�S��fKگV��ގ��yk����銀޷d,' ���!�
m�37�^�4�1��8;��]rfd�:̌X2�bo	u�H����E�C ����&�2�2�W�uE�J]��\i)I�av�|=#�Z���ݬF���1��Vxh8��{�l������ޘ���������p�����f��_�l�� ���znl���A��C�2&�V���7+��!����f���9\��M{����-����>D�"��[=Ku�@5�i�H���7�8L����:�۶0���/.��3:���fޓ�T�D��b�e��[���~\��S����%@�����͔!"����G%����$z�)bw&�v��'ۆ��7�i	�M�T���"����c��jD������LF�F��
�!�4�[t���͐�wFd�o�T6��s���~���f�Q�I�s�����M�
L	i�G�Gٿ�T��'��ʴ��~r��ƟLw\�)����\uN�@���G���M�s���	�̥�M������[M	]\Y��U��d�2�a��$qv�� �<ǁݑ��
hV�o��(H#^X�@T�d��kl��ZW\G���\�D���Q�>6
Ѣe|ǈ�R|Ȃiߓ�_�Y]>�h/��I.��ՙ>�p�g%�-�5 ����g_���&Uӿ�4�(�zs�A؄���ɉ�Vpj�E1���x3�p%1����鈯��vBʅ��F&U(\w��|6a��IhDI|��[�1Z��D��i��q��}]��ߝ,�T�y���ݾy�*�7�*��n�F@�������<���ε�*�22��$~��T��h�s�&]E�Vo(������{}��
��o_H��.O�] k����DhF?�n�YRq8�(vn����0?����`��ƅ�"o�̥��cx���E�Z]���l����@.dd�)M�c���D�L�k/�\�>"Qa��K?6|��q����ff�i�y��XC���Ijq���>�Sg~��hr����ř�N�f٫	ܛ�ݲ��~�1�#��p$�yؾȵ�s�����d5q�=�,���t���iyN��Nj��tL�/�ﶵ���ɉ�e'�����vn�,�·�_Y��s|���~���t���{n0�c�����ŢR:����݂w<L��*�i��\��t~'�>Y��f�aPꔴ^*Uk!��|4�����@�v��A?G
h �����ͣ51���/x�3�I��h�_����7�*V+t��]����F�v�:OLM�}e�$�����Fv.�͒�O�R�<���u�F��㖩��?���h�6.��"���vkR��5�JYhh�5E�W�6Z^���[��)�	�_~���3CB=��9�(5���������� ]<g���������v��8U˕�Ӵ��{�nӺ��o}���
�o5��a���� 2�]�E���5P��cl�n���S�6_!V�}�#��bi�j�h��Vԋ�Qo��8�0㓲��._n���7��aD����C��1���ɱfM7n��k��;].j�k���#2 4q��7ȃ�̝2gM���%�G}3o�C&³j���b����I�Jb�MkZ�i ~ g�>e(�����������ҙ�7/C�Yd�~Z(5�7Ii醆D�*�A����]��X%9�E�Q���w�[�q�WST�A%+�-��/t�b��I��������^�8��X���L�{���EX����`�>�1Y��$���? 8�M��gP�����{�#���"/h���NYn����7�W�$hu�z�KN�B��N��� Ѐ��,l���f�b����gkV��5ӟ4���O�pG��ø��s#�����>����.w|��Q�LBR7:���O�Mݽ)]o������k���s"�ΰ|1:��f2O^�����H4u�zGN_���p�����Z�^�?�x�b��������v��`�<�h]$�89��o����sf�
��2|�S�zE�����e$/p���`��g	�s�0R�ĳ�{q��Ӡ���,NA�����ޯ֓e.uǹ��*����{���_K���qG	�2���eT#��|��Q��N� �3��C�Ņ����[S���hi*��8��L�
e��R���T����sV��3����j�$m�`g�Veۺ��v�R?�<����C[�5x%���`ۊ�pq���"ph����in�/'�t����{0>�����AZ�V���L� d+�4eO��lԨ#��^"��܏�ZK�7�G4�����.5x�Ά5��b}ꁋE��`ShQgͨ���-j�&��v�`VC�+���J��z��9���"�� h��F��Ӷ��D)亢�3�q�$<݀�5D�x!"w
>��+�.�H;�h��/�����{oCۺ-U�縯�q]XX��Rk ����k�ފ�������D �`���.�x����m�%��x	��>�["���y�ǲ��LW*�I4���I��!��)f�� ��G�m@ze	��(ح)��tX��n�cNy��Ǎ4]�?��sH��E �#V��t�Jr��z�/b	b��c�B��;��w���$s=�~s��*U��Sc�����!i�5�����2�;���^.ߏP�Nz�yE��ゞ��=[�9$��y+�y>}7,�mw@^ͼg�����~{����������>xT�ݺ��#15��1�߃K$cv�"�q��O���zn�~�������v�/b}�3H{��]�N%�{5�}������4'ec�L�H+�8�����!u*���)��_�NM6[`!-c�FW_ 
>wH�n>��Xƴ�j��3A&<��CI�G����7 
��D�+:��~�p� �=���,���={��[����0�%N�|���Jj�O< �I�\'V<r��(�p�z���&~��S�e��N���*�xo�*�ǉ�wg5� {�ۏ�'�|�d�.�sc�q�Ƿl�����j���EAT�D���R�w��+H�5� *ED@A@z�%�BT��tBh��Jh���A�s�c�W�=��R�^k�������=�,��jG�Sen��S �ۻ,�K��3�N��|N�!|,�|$�ΜcB�褎wI�7�i�$E/(	��q���������U/����l��mM�˕i���r�)�H!����]ߡ,�-R�P�{�{��{��k�ec�d�4:���Z�~��?����G� �0�Re���d�
߬�SE�#��G��L�X�W��3y��Nڒ^�P&؞y��/D�L]W��ȣn�>H֦���aF񎩯/qB�	h�:�?K���U�O�g���.�nkH�����³�;*�2�3��a�!��G�`8e�5�)�-��q�������u#
��I��`�y�:����t�)Q!��S��N���k�5Ғ=Y]%>r�F����=�q�\��l��h Z����% ��@�I�]���!����	��"���!�6�@ڵ��@w���7�_�C:�M�&��-KFPf�1��!�n� =�A�ۋ�ҋ��Wyy��ӛ�p����5��I��8 ����!�D�����[Op������\���S��P��@���k_zE��I�n~�1]��lI*L~� ���R������BZ�x���p��>v�&�����ʒ���R��K��-�~�D�b�� '�<9��?��E��:'�o�����}��H�N�C�>}{J�F�iL��9��  p�Z�G���^m�J6�ӏ�e����؊�zb�4_�2������G*�.s�����}��0إ@�$��;����*ʎ<&d�g����[Q �lK��'^b�Wb�h�n0]�<�����e4���O{�:�^���I�J��5X�M@�GV��}��G��c����Z�����ѝ�N��BZ����B�	�|�R(q+z+��F+}ނ�M�jaQ�d��U�|^��g?���6��z��Y���מ�M��<�� 1h[��xu����e`����)BH�$��٘F�r1n���)/�=�qu%XC�+^2߭�R��v3K�1Cu>�=��J;Mͻ��Q����ܹ=��)Q�\�!v���SE�ξ#�gs����R�T�k��}-�i�3_�n7��)T��B�2���=N�뒼���Pza]v�m��ۛx%������/�o_�Rpd��X�ʞs{��@B��ok���N�:�J�}����Cx&�|��5J�qN�) 4�P�W�����[@��(�>WD(jd��.�)t$���Y��T��3�)%|��b������
�>MFq�=U�>~wŤ���1�\AZ(B���_�O
��x����ܰ�i�WPT��n�s�ܴ��#n�Q����!�n��۩xܔ�%�gT��Ǘ��s���H-ҫ�Tgʲ>.O����Q�a���VC=x�{�T�5�jc\��ٍ��X�-
��-[N�6x�ΕbeHvs����A��8-���	e�k����f	����\cD���P�*�:�=.fT�޺k!m�
�F��-l}�W��~��	���Y��#[�ߏ<b���ŉ/	�Emmԛ��&���ў��eԨ|��)�r�_�A��b�a�-RSkH(�	�GB�cas1�A;���U~�0���utr?�\^lK'�`C��wi�\�&���{�dAc��*S?�9����f�w��,J����^>:��,l!�8yC��<w=������))3zњ��:�l�s��:0��ycm��cB�5|����<���7k���b�ל؂�.RK}�?}�]V�����kr�����9��}���d�TT0\��x5�k�g��c2I�ӽۋKK��gU?������\Ն������*�Ŏ^��r$�zq
7vt�UyoF#�RR�wM����I����{��A�C���h��a�J�[��":e�����=8���T���?8��2%���������'r�ˋf�BZ3��BZY�h}�|
��&8�>S�.�o�ͻ���O��'������m}5�c�;X3���m�zb��9J��2R��o�����|% d�xq���_^��y������{��^�'ĿxBxI�⛇2���H�L/>���#y�����jh�~���%�z�i��$�j+�'�פi��c����N�io2j��yCM�y�)&A��|�U���U�~RH�cF�����=$U��A�����$	�����!�ǏWu5�_D�{��F��Ab�8�t����1�1�]�������s�2N����J&�B����'��4-e�*~~�וh4dF�k8SV�֖.oe��~$���v$T��O�/�R��뵠��gМ�:t�JE�Kŏ�c=�&E��i�LaZJJ�������~~Mj�"Y�)Bʱk#%�D$�?+���PX	"I���O��L���&��&�˙6V���1�k���_RR������������G?����=9�cb���ϰ�������y`���ڴL�~�q���}��Xf\mԸ�Sk�����  ���`z積1�=i��^��,,}�Si\�OĬ%RhR�t0�������w$���6J��PEͧ����'����V������X�ii���҇z�'��nP\����*�����3�����Cf�����9�S����k�����;݂�P-���4��O�'8R���Ƿtgc��ua~s�zo�^�ώ���djr%���au�gm�O�jZx`�^�˼����^��n�TD%Eȱp����g��(ی	+/���܄�h�m}��<�J�K����0�d�{L^vo��|؃�6d6�F��ϣ�����N=��ᾒ�;�F�$'����*�ǹ�a�G�5*
� �&�^i�Y���;9�>����4� �t������U	�G���/J��P���b�?��΍'�^�lPT���xM'{�?�ka����%�{.S�'[E��Z��ۛ�cy+L��ʵ�2��y�Q��ڇI�ݶzm���B��Q�Mo�X��՞�Rl����%竤b��;����0�%���	���;�̝�Ȗ~�e&���/���L|�^h'��ш�q�y�3|�1�  iX�z��\; L1 �e�̩ķ���71��qx��C&��_�,��wML����'���k?��ܨ�zb��J�C�p�C�|��#��>�8o�l�d��P�YF��wMsҞ=��h4!є�bY��棯�^X2�'m���a��dK�n�NJկO��t��ĝ�QKL��t���+��#�����"�7��\�L��%�� ��J=d��	�޽�@����Dp��14��B�>����_"�DMnWҋ�*���@���k��N&#�ʈ[�ѿxp>]��f2�)���DY}e�3��2)zQ��x"Ϟ����&@>խ^*�]L�TPX�ſ���~�w��łR�Wo���'�v�%�=�)b�׬ H���8����Q��j�"�;
�a]���nP\bb�EL��:WȲ\6Xy�f�T�"c���{�/
���������g�=b-YZ��ؓUX.��>��T��U:!��x�f9���DHL��6��)����Ʈ�:"����F.%jp�IG�d��R�&����a\z%�~e�u-�!����)�7�Xa�JGW$����e�P��&�FGǎ^��,+�R*$��Fo� �~�	f��J���<~�M�vd{E�իW�7���Ĝ�솬w���D\�1$T�	�L?~��)J�F{�1~��O�Z+T��j&�@yR��ro�G��臥�J�d
�j�ڗ��L�NTք���0 |�Z��H>���=P�"-����\*�U�k����;����N*6�P]d��ؙ�c�Qd�`�9;� �[�Q�֐u��S��O;%N�5�B�+[��Qʤ�� ��}\�yU�����s����Z�ms���cx���"g��3
O��t8'����@x���
y5��v��g2��Z��s�A�+z=��`�6�Jۮ(������I~��%H����>�/u(��Ih��ܴ)���>E���r��7�f�7�M4��3D4%�����5���)錬�L��?*���u-��q�"/�oF�v�<ο���\���Ԩ{8�E�����)&��*K;�����@�l�)���_�6��܌p?���.�H��0�}o_�'�������Pɋ�����j}$,ژ��_����n���G.Zݽ�&�s^X�ouР��855U9jy~=�F�yV�b��z��տ���zl�a����1k�[��k�ɩq\��U��߼�R�9?��df%�����5��uf�իWB�➞�x���#<k8���8e%%=�0����p4Z�:�B{�5?l���$'�[�&j��;��!i?��^���H$M��p	����A*T�â҈Q�mT�z|��GpW��L%����N�y'��͚'Tu���oJo��)�=:�C���Lׇ���M���,>4����~!����٨r@�@����|��}��?3=r�����/�����dYe�|�ʓ��C�O��	��������Ǡ����6�vj��㗷�5�{��Ւ؋�I-#L2A�ɡyMPr�gFщ��Pr���ʶ�ӂ�d��������?�N�!W��""��x�O �^&���|�v�J<�u�l�r��F9C��#����g|�M�۵�#�:��M����/���|d�����LÌ�|o�krW�w���z��>�:\����Nx;�TV�8�@<~�,�y|o?v�GF��������U����'�ċ]�Q���>3� 3���7�@�o��̟���D��Eb��ŕ7g��>D���@@P��X����E��`�V����ʛ6������63����C�7�cf@C�jt2՝#p��X ��x7ٳ~c7��1��W?��r16ˆ���3o�?�m�ZKL��*�����U��{ITm1b+����k���]|���Sp�� ��~�9�ؾ\�׌g0�������;�%����	g�UE��f�X��7��}�k`8��z%��ǧ�����r�rm���ݹ�oy��/�V+8�G�F}-7�0��~�;� ߯�V|a��4�+�z����X��M�'�c d|��[8�M�/��2�� Zெ���RN���Cq�!�/�<=Q4���.d�qOqv��+�>�_���>��R>�D~�$���1�GE,h��MP�����O��wl1���Z�3�i�� � f������V����y�?z�Z�U��\h��т�r�f7e�������u���q�[�5���O	W^^��a-�X�V�A*?�^q$.&F�3n�Vl-����d���#Q6�N��1�he�g�7�ǅQO�q���NЀ8��Y�;���69�n��z�ZQ>���!́G:^/���5�J�~nz��H|f3�mw޴��dSP|zc���KZ��m/����V����C��Z��A�b@@3	e���7"NɎ�J�˅��5�:�f_��߹Ɲ��5�w|��Jf�bW'Y�9ب�'�εz'����PΏ�z�d��74YM�*�:�܋�GG��"��+��mx2{��P�\̤�&H�4�"KS=�Ye�;�CIE6��ƴ���ҵ(D��C��H��JM+�e��:��+xݦX��9OL����"-f��@gBO?P�$����o0��"���������u���-)��wPi�ym�OТ���E%�Oa�p`A8>��	A�	~��7��P(�N�W�A�z�71�=��`6X�w2�f�BO��*	���Ϩֻ���]y#%.� ���VH�g��>,�|,V�uU� �[���P�_�eL�_��Cv^�h>�&z+��C#o)&�\[:o�3�6յ[XR����7:�5�=�ES��'�?[��`�Y���ܻ/����������g6 �52zL���^[��i�SW _�ݞ�O<���32?�8�p�&��D�&�щ�|j�scrv{@������QL���y�@Cu��G����ϿJ�/���o�)o�Y����>r����d���9�1�>�v��� j�����'�1�I��B3��Z;�?��@���m\�>����~J���%S1$���H3O���Z���#r�j��5*
��� w����V�.@�m����HVO����s�'�x��y{���=^r��Gj�U�G�"��}��Vv_I
�B��T�iv�����V�kQ��l�?E��i�[��QM0"�����1��̬�{3ѧ�\OaI�dl�$J�0��k���'B�a�' 4��))�)���]�X�)��w�߲��ON�|�@��?��Ly8C$IM�T�c1x|�3 �K5Q/[��N�����{��<v�%�uq�]]�o�܀���++�q�~$\~#!)����cO���홠�m)ҧҝWؿf�"B��6k��P��րχ�1��Wi͟�o]����-� ^ׂ=HT�2���^Ȗ�U������˼��ݰ�-.|l�=/�(59z�oJ���pY�ބ��������o]�(ص'3��ֺ����}�IB�RJ�Ѣ���52`zhH�TL�H��~�A�d��4�+t��+ی	XմT���B���[��\���cn�+u��mqwW��R���.��M�zg��4� �E��'�����l��Mtm~P�G�+����v���L��=�a}[����	SN���c�/��#�ӊ�y9����[-^�'�B�c�rNVc����xM[��%��!���.�7��3S���ӥtr	�����&#��=>VK\%���T����ƞ�w���W핖�E���P`�zHUȗ��!qK�C�(f7�Х߮+���9�a{?�B.��Т�@ѐ����U�2����uv*n�T���gJ��)��,�Σ�3,׸�2��;�ds�V�_>����`J�������w�7�j�e���>,�z�����+���N��4�(�z��I]f�S ������r�ʽ	쉶�i��]�i�댲�����rϙo�=�m�e�&#h���|�|�$�B}u&K�� ��٧B�뽖��'9u���ڕ#��s��r���]ɓ�����>"j�NQQS���Ŗ'K�V澷���tI�kv|�(>C������%$'��Sꞡ����J󐇛�z�N�	Ʊ�<K�ڼs����3N�'v������ַ����^�Y i�����H�`�����G�b�k:�:��}����\�"@�]�z�iM1�mH4��3�!��,k�Ԉ����b�_ִ��+�<7?�XCtޤ�ω0�5.��l"x�F��C�C���Lm�X̢���2w�8���i��^��>֬a6z-b�R8��d�gZ��Z��z���Q�jH��5���v8镳2ښj��֋RR�M����ץ��J�yp¶�{֮�^�b �.���7 ���O=�t����D��F��5b0G�$���y|�ܠ.-��U}����Y�[¨G��Y�bHz��K��f?M5�Y\��K��f'�������j�q p��C��H��v��K��j�6�Q��C�f��qP��Sm�d,�.�:ʘXs�F ���;�ؒ��ҽt��L�����)�M���6[��h�ëۿ���,\��c_��l.<�?�N�<��̃Tb�1�ǒ����ɂ�q1/���J䱇��tͻ�{�>c��Xr�X$˝ӌo7/on	�7[�� ߫����x��8�@��ZѷOƸ'�l7��`vR��G�P�5@f@��2�D�'6��X0�m�"O���R=Ǿe��R>:i�5�|\�r�%C���LY���y����m�-S[�V^e�*s-���_�j�f�Dآ8{B�˶���T��ĪϷZZO��k����]��M��*��� �wl��nc����5�JO������$����6�(�M+z�҂V�";���Ϡ��W�p/�d�?/�R
��ʿ��^�pH��+��*���5zd6K�	��iRe8�$l�Y�pD�O��"p#�|��CA����#T��1�C�)V��(1��Z7�upߙe��Ρ
Ł��1�o�shP����p�Gkmkjzm�z�����6��V�������5��:�3��j0���G!�1�����Ă����>�����V��������BN���K�C9�F�CS��j'�YD�����=U��z�*�o��f���.�[B�9L�~�#7�#���:�ܽu��Sr)���go���w���h�v�V�)xsʿfr�P���u�#O��v��5(��G�4~[ЪK�҄�T��xu�E�wWM��|6�R fs��)"�E�c�֏���_�Y[/�4&�|)ryef�޴��L�=d�`��A��=X�b�M6�W'>�n�>j64���P��@}�L��&��!�%t���
�}�����_C�Nq��q]G�T�G���{f��l	�b"��jc�Z籟�R'6��&|���>)*�zJ=��p/Ȩ�7���fKve���L�"�r������<.�Z{��ؑ�IR���A���>l��������6�% �r'����6�F�Lw�gm��<8=SQT�ez��\���QY���u/�Y�>;^��\Y��<�Vd^������4��*@�<u�4�[��	��U�1Z�pĺ��b�N)2uXF�]3e��Hm��=(��V/�f�n-ߔ��������n��6��:�r:����]ss�ޯ�o\m�'"OM{{�U��#����~!���t��%#�>�&�涘 �"��%�ٞ�������IZW�o@�_���XԹ�x� �1	�׹�ܼ��!���N; �*��A�>�j�B�<�9zۦ����+ut�>ɘ
۽o�-��q�����*�Dŷ�b��@+��)��K��y�[�/GQ׈WRS���x#�Ej��Z��㏻�����r��]Ex"#�"*�S�N�-�Ddk��g�#j�Ï��P���s���\�-���˴'ּ��tЇk/0���6�U��eA��>�s���?�9*�ϡ���;rh�.jz�{n���,�#�|��l�c5	A�o�
������67���e������7�p�	Uz�2;��I���,Y�=\WO�YEc�ײ�ȥ�C'4��X(��f��k�dT�E)��:r�i�nX�V��^�s�Q�����Hl=q�wz=Qk�t�
�z�P>�EA���:+�U��a�о�}��ﰠ���-�@$�����\��<9��%�$�s
��+���P��,�R�ʝ2\��0�}�J�f��Ipꨣ7��x�@�؉Y�������g�o߰��ի�S��hV��Y��=bZ�{�i�t�&F�K�/�u���t�3&��\b����V���W�fN8z�$C������#~͓�\��

O�~���<E/]	DY��P�<���d8i�H�|E���m��-A6唦Ӻz�^w��y0.��@�~��5h�`�@���VՍ��/�/6R博�����y׋x��#�3 ��͌���Vz�����#�}���4;�!c�R�TD)�.����	��-aL�g�^= "�y[��I	�Ҝy(+�z����d�Cl{Ֆ�F(�/_�7;r4M���$$��3h���1��L<u˧(t�oe@��a���ٝ��MZ�F��A�
ݗ�{�R�W�X}Ƙg�j��R�u��k�1M�A�ޯ�0_?Øz!1c�V�"���v)��?z0������oЀ?l00���'R�mҔ5H[���*`�~��>lv4G�1q�7L�叙(v����3_�o���u|��?~t,ț}C_, �sG핻��g\,ʎ��s�ؗ�8��p�r��&o��2/�u��'���o�q�T:zY��f�_��c���kN�V(��ijT�5��'�"4 Q��*���\�l�B�y6�^��#EV�H¯j�����g�Y՞���U��;����\��<�����]'q����yĩ����݌gsq�(�`�J���qM�MI,�h�N�ؗnD�Y�ln^��(�i�����PBXX݃\���b9����I��ӫ|$׶K&�3�\ba����#e*��7Vk*-5m2 +��}����fc>����U*f`6Y�"����)��6�Z
툅ו��/T0�0��>G:	z7h08%�Զ�)?�r���{�S	j��LM� 4?HW���`_h�s��I@��Qs���i1sk�Y�Y&\��}���2 ��(�pRDl�܋�d��r@6E�)���7!d����r�S#x<N��.ܽJ����0٨���j�-8]mt�(�Th�Nbn������~���}vP��-����%�Y�%]�� ��tg#�ܥ�-���Q	.բi��>߫���Z�h�d� vW�y"nrʱ��g��x�ku���X��a��%��Ӄ���%�ЁXTV ƇP�U�Z���3��h��얃�����f5��	_�E�V�t2�P{�^�v)��X�?ȷ=�r
뫷[,@ Y�; �T���޴Gդ%��Ѐ�;qУ Z�+ܓ}4J6vP.;9LAS#.S%��[����ljA�j�y��q]D�)�k]U�������79����|`���J:��}n�r��.ט��[L��CĆc�Fu�;�+f���"��aX�^�� �+��̩ʻ�'�� �g�8�4f�y˶�t�?�c�|�.i��(r�
��d6Y�܂�]��S)!���[d��M����p�ʖN=K7�Y
�8W+�n��%yLz��:�ϝ�����I�(��Z�$= ��k����m�q����X�1��r��ͨ����,���q�?��ȓǜ	Ks�|� Y����8��\Ir���U��J�3$�YЬ��$����('^����o�(�K�I]����x9��-��-&�e�J��[�������J�))���Z�0�+P�}��.��f@-���Gg��"�^HdVk��Y�|X�f��$k� �i;�Mk��OGj �9��ǋ Ӌ�%|i�\�UW$�?Yt����aZ�>�4p̕x�f�asҜ+��|t|)M�[B�q���o�|�Sļ��T/2�j�\}*���`RO/J�f%1���͛@��;�8����*����Ý=��wg�u�s1����f��Aɢ�n���.�IO����@����e�i3�e�ZX�����,,����%�cҦ�<��Hhn�In�d9�6`�z#�؂%�'È�-�F�7��ʫ/:��@��q�)�8/Ib�-(��:�J��_�o����K�#�!�uJ/��A`��vvIj��S���%�+Uc~Evj��d��c��ꌵ��>�t��2�����`����<Q0����`j�{|l�����zba]�E��!�:=�νSdKy�o�/:,�Ald 9�돦ٸnG��;k�� ��l���P���t��$����y!r�KƐb�yi�5���ю"��	a0�p8�u�ԡ���p���T�0��#�'��
��<K1=9��/<MJ��/\��^ �����OYn��o�����"v���[����Y���ef�\�u�}�l�A12�i�.-�t�g#B,ފ�pOdn%�ؓ�"u?������k��a�1���B�*�+���ð���
au�Y��|��w�5Tu��T]f�}�Jº�- ��N��L���/Tz�њk�^���O�{�%e���p�S)BH;% �<ۭ`5�B�S ����Q������mx�^ǉ�����E�3���F5�*�C}r����bC"�Zs'lȁq�LC/['��?+�u�0���Xn�:?�u���զ�Y�S\N'���e�2�Yv���F��n><^}���O3�Z��]��	���+'}�G�5��{p3>�Z�&{g�Z���|���mJ��^/�p;5!�
%�}�g�`�"�7��HgkÃ�D��Zk=��Zh}��OO�˫NL|T�뿙���������8y��+��.����k����u��AK�ˮw���B�3�t�y&�����8n����ϛ�U�&�����ǢN:��%xN	�n�%Í �1VӬ\�� Q_9������U�O�m_NGӏ�[�vB��mJ�^��@Ң�K�X�1����!��O�B�S���"P4��Z�O�Vf��R��{���*����ߢф�
�==���F��&j��;7X���#3�S���UK����gS��%yf��$CѦ�7����������\ � �W����ޙ�������A���c��T��z���_�vK��]ݐ���:��n����Y�(���k����sJ�rͲ�����t��j*MJ\\��[����׸�^�.|��
��6xic�����p�#kp����][�V�H|�^��]qau��R�-��nUWO�P5o�#o�zm�.P���Y�Թgz�Ɏ�j�_a�Z1��׽����u@v�@��������H��ck��W.~;K+Y�/�l��3]jg�=�S$2�D�:��+�I'[����H��S1@�ѱ�k#�y���7A� �@kbN�6��:���ϫI�F(��{K�q�ڵ��)vI�6>�<�%�?�'=�cz��܌�p 1�<c����l�K����L�Abꑁc�'[w
��5q�D�)�E(U��像�[3p��|b&�~'�r�GQ�g�{O_4��ċ��f��P䰿IS��W��ȱ{M�Cʟ~D3K�0�)ּ{ȍ��,:�'���g�Y�rzR��ԇ�6┍8�A���z���:����mJ�&����Zʺ�B~۪���=L:<*I�z "0�"g���oO�~-ɥfw�csQ3�DhOʰ>��KGX�`��P���ZY��m>re�lÏgD4�7,����0oee�Z޹Mw�2�q�,N#4���6�3+�����O;���1(���)��~v�C�UL�Cj��gN>�ݾ��}w��)y^���QD��L��s����D�z��	�������rS|m�flC��_9�B]�+��Y���&���+r��&8��ϫ�}q�q��Ag��a��3�⛱Z(S�����r��p�9e�|M`�@;`�?����B�Dg�w.�A2�d�,'�J	�e�D*��wbT*45��z�`�C�{ WSRЉ1k�b�#��zN֨j�g�R�ȮR� X��=5�ed�;� �n�?:����=x+�AU�h���ˤ?���a6��7�*���!o�lv0�ۧ
0�)V{�xn����%���?�.xbtӛ� 
%.}sAN��k�!������p^^���Į��EYC���j���R�7Z<?��:���QK#3��-c���}Ѐ�rM%6ȑk�� 7M�����0HR�`(�[�"�#���-�Ε%5������YU�K<��n���,ֳ�|zp�\X�����6��jOj��R_�/$X� ����eA�D'//<���$��l�#��ݳ����C��A�C#D�������?�qD[�A�����xK��k��1�O�է�̲��Ջ�}އQ�e.Q:�HJ�Lx�|`������oT%{��C˴>����%���6�Ꞇ<eY/μK@����o�&ce������X��i�,	m��k��}^�h1s�K�n�>��М�I�]k>_�$���y��&Zp�;��#�v�o�+�����p��0�`�=B����������qH]RK]��_>O@]��Y�֦M�ȱEN�r<qi�:��Z i Q6��lX�%`;np(j�3�M�����/ii% ����il�Z��b9��8�f=�4hD�����<���:����Ma���!a��W��(�л��gV&NEs�ΏZg���Ż�|�˃�шj<�:�U��1I�aH�퟿,���Ԏ���"��N��w�?���\�h�y`��Lf#��m�*�Q�^��ngq8K4/��������t���;���
��X>Q��h��JZ@&�y@ܯ������ӆ@�H\\���%'6���5'������)�D$1����!�v����=�IH�D�h���҃����B��q�B;rQR�H��=c��EƤDdo�Hz�.Q����\�A��N�[{�¯i�۞�;��(���E��f}��vL�^� �0$���!�z$ �O!�Օʫ�T�,
�Y
C^��wۀ���O� ^�e�e��b��/���m���l�l��μQ�L�e��Ņ�ZS�ev��Zq=���nR���x���ݭ}�,����� '�R���CUPb�ã�X��5�ئ7���]�ρ��m#=0s���`�������������s) �o�K 2��}P���� &i:�����j�p��(�媆m��m�^���̃�O�b(OB!�3�qV�] ��.*�� :����G|n	����h�I{ɻkn(��5�mr��i�v�����W`��,��cR�>*�k�'G�ڀ{��w1�r�kʟB3�s=��*w����� d���������
�t�y;mh����d]��ٸ��������-Q�M�Q1WH	�A�x����;�#E,�eDD��5��z��rVX�������B��ܛ'�'����w��V���}*�:io#֕���Z�A&���c�LV������}������.;�/С��K�}�Tr�8�.��7��M�L��(����'�vC|��#}T%�J��9a��H�%��{忥Z�Ԉ�Ă���c��ּ�[����	�`�Õ��rb`�^�4m5���&:�^���������7?�76�%G�[�m���i\h����X/0�E�Ը��D���y̩�ܻ�J�3:�2#�> ��Y���Z���j;DW����7�q��-��N�'c]x 8
��a:X !�(K�{̀,U�K9|ZI�$��O���8)��"��0�o��po~���c>$���E�H�����-p��^w���~{A�#N����ö���󢉭&&q/�����<�Q��u����C6���*HM�:��T��]Zx�<�h>���1F��`)��T�ڋ�Y�o�^|�u�I��<��ܰ�D^d�@>����c!�ί����r���Y:��cʒ��{�˔�=D��X�������T�[}�R=�" ^���bV�Y��~Xm����RD�0G��O���ަ�9�� �i��ვ�@׉S�n<���N������҄���/�U�ИD�NiȌ�}d�Ɋ_|,��1UL��@tF;'.��_��涴��8(Vz֭׊8u�<ꨅ�댙�Xq<n��Z�[0�XX؜�c��<8��V�c���w�*�R�@���2���~" _�
l8 ���_�%h�c �Hu��K����LL��
x��L��9�>?G]�xϒ��^X�X�B��W[<yF��	��*���I�����pߡW��Q��i�@���#�h��3��~�8�����P�jP���1ſg���Ʀ�򫝾%V�G���$�-��sӬOM7�p�q�����jL��>��AY
��?��z��"H����(on��#�|'���c	3��bL|�4ڬ>?�5S�eQ4��UTT�A��~��l��w]�z��'��mʈ]#��!~p�L�a�,��+�س��kޒ����V&�ꟀGiL�*�{拈�a�?���F�l�c�2��敟J����[��>:<�iR�&�P��e����4���99����&�0��}����������t�º�����T�Uʆ�MK�${u�Ø��@`�1�{J��U�&Z��٧�-�V�.ϳ��~���A����LNJ���M�M�X�1W�V�x�����k�Ap�có"u~��u��@7�M�,������j� }������s���=�Ԣ�28�#f� ��������J�9x�@�ğ��P�[���\�3i��hqr�2��wx���l~l�*KV�{���c/��,��F_�4�\�ތ.0�,��U����8%��I6�^��U��>�|�G��r����S�l�N�x���Fh��|�1p�*��X^�s�Q񊕈�=����	����\b!c[�����{���XU��2��v[�65�Y,����z|M�у��������`��p]���p�=�\!v�7��<"�C��}�<��ܐ�v�X�:���s��;���4�33�z�Չ�_�B�����=8<�1�}����6@���Y��x� �D-K��3����ދ���˵��Q����"`������ƣ�!��LK�C���{"O�m�҇���j��	x]�~wI�F���O�|�wן]�|!����+v����$ro��5��/���]
yCr{`���Y�I��9�˳��W^����0���|��2�o9�	�����D�B���T���7��iK_�t#�Kt��1{n�-E�O�Au9h���,W7/y��'�/=�����;�֋fB��u�,Ά�v�8��0Jy�T��ޅx|������'�q���r�IM����������*��t����}C	��I�H��[�~?���3њ��Q�Y�'�<��� �v�:go��W+��V�¸�<[JyZϥ���_Y�H�m�|fq9�b�0]�9Cȗ@�rUk��wi��U��SPý�����'�蛥=�;�B�		��x(��}	)�W���u��]�F��Y�k4���V|fu�}|5�ה�y3�sk�B������ ����0>���Ծ�v"a�󷫼��.-����f�]�u�C�����?�tS�
_����[�Y/G&�Yq����cPa�TA2�Ǫ�����ڕ��?�|���jT���.p�0弛5�P���q�9�[o�N̟��(Έ����~����=��3^���ꭙ�.�АKb"�T���a��w�����Ņ%;�\�LYB��"L�i��L潧Z�o�2o��8��|�*�ǁ�����n{d��&����}VV"����*�"j���+�����>�$XZV��s�?�96>��ߗ�2Um��]�:�,�%����������z�����c�/"*����+�:��(�� ���w柽�����y�tu��%��������v�����
�X���tp�[�'����7������n��:�PO���}+������x����Ľ�2��>�ۖ�ou!c�v�����{�!|�������M6�q�������Tj�Ԥg�Gm�������j�އ������CBZB��������K����n�z������l�>g�Z�z�}�g7Hg.��ұi�ӐHd���م}���=c�ՋE~�),ȫ]�-�W�u�NN��u��"8�h
��y}@���G�������X����IXO��JSF \�8�o��Jr,���O����0��U(�@��y��^s�T.�s�n��/S1�Svھ,gsqÛ�y{6��� ;�r���������c������X3�9��s��'�p�1p����36:��9:�F~n�jd���*�qWo&��nWp��]��S�+3��L��	�=|��]�>�-��M��]o�~Y�U�\2��)G����"��`���d��=�`oc����+Wc��O`|�<o��U'�!�� ��c}a��\�(��,3�g+h=���ɨ�L�I�w���(�k2�A��(b�FEj"�&T݌����c���F�ᱣ�cC��+K��4#�� b0nK#65���Ǝ����z���Ȟ�0����o^5獽C#,�¶�bP?	�j�R6����Ց�s�ҟ��4ᒐ�D��CJ*Xo�k����%�<$��Ƹ��+��(O�s�j6$�U�F>��.A�\s{�7%��yy�(�)l�=�B�=���=���y{�e-AxrG0�Q�����k�*��a^�]��f{��砗�ܪ~H_j�l����lg%7��oʠN�����]��~�zywhs�*F7�:��wh�����d� �ϥp���Dk�5w�I���N��N��N`�\�n/�,�-V�P��6�42���&���o;�	�GY��t;�y8#K�8�	�a���.��&ێ�_��<�ir�׊]��;��\!3��z�l���ptG��)rI��֢A
�
~g��VBn�B�F:�L?�/93�$;�����dN���@ܿ'G�5��7c�=Mln��g�Gw��Ǽ�����M^����S���ɴ$�+i<.x�C��u{��:p6� BC]��LBFBY���pa����y{ȅԿM�]5����[Ն�M�������4�#g���X�U�fg-ߞjܞ�8[/�A��D�樉�$l�̐ۈ�m���r�~�����������6�nd�/u�z��߫Ȍ��6?�
A�['4��D'���e\�l�:`��܂�����Dl����|~p������D��[�l퀻rff]�ן
l-���s�`*�����uM���2��I'��$R	C`��d������֣7�_*`@�6GQ�e�!i4'_6��(d�֓96��;H���S��N.] $�	2'�@��4�18O�W�n��T�	0}XNB0_��@��]0�Id�n�`-�o0�`Q���+��J��U<<<��)H�Ŕ�uY[��fw�}��������R�Ep�D��).��}���,+)=D ��v>�b
m,�p�'kp&h�-�4�0G����S�hmW����>��]U�wb�eb�����K�Vפ���{��Z��ͼC^�H��"i�}�$�;t[Zc�u���<˨���ͣ�Tkzkw���'�{!D�-�ďS�ꪂ9��D{t����o�9�̊IΤ���[Xj��Nv�d����x�۷�]�ɷ�	L��K��GX߶�¢��r�M
��[@tM�,"�-��a۵?�!�R��Hd�yو�:WO��8[��0�/S���ъ�,�dE��T�*���YBrYllB�h�./o���Kt���ۣ�-���T9x���'~��i��:e�K,� `�0��0�tȞ7=��m�vo~����O��,쁙QUkc&�S��E��������=YHR�
���g�n�lgoP�w�[�@�ɲ�B�������Ê�%�(��6��=�k��jg�V�l��K����JY�H�{�pp���C���2�"m��a�?w>i�xq��D� �u�'UB���ձ�L)�|�W�Qgs+��+Ԛ�L7M�ə�yD��,��/-�fy��O�|��d5#[3h�D:��U������	��+m�@,(�ѫ�?q�O��y���E�30/ �������BWS�Kq�#�07fhfUQ[Aǟ빧��7Z=��Y~U����IԷgaA�x��w�9=���-��w���FD ·2��4��so����)B5�R����	�'�cӉk����3�<p-��|k�=_x#�Վ��7��Tٳ����j����o�ShT���@_$B���|�06&����Y���#���>	�t���0���n��>���O�6�Wa�0�-T<
�(��}gg�ӵ�C������H�%|��j�ɿW�P{���N��o�ה�<�;��u�}_�j�]]���{�:��l��ν���F�׮�ec>���mӢ�O"gy5K>�}�`�|L��	��0�s^q����^^K��LY����Zyj�]|�O�^�w��v1q��'k���y�Qo�v�s�n+K��МI� �DQugd�F�����"��oBh�9�M���UR;�j2.kԷ8E�;p#ր]�.T�j0��E ���}Y��'[�Q��P���A?�G%P���c!�{`�nwP��1�&���{t׈����)��E�/O^֏`�?&�>7M�ea�y���J?6\��[�e�2�,�H ��5�;]�����/_6�,��ڮ)J}���*'6��س���N>�����0%Lz4ʙW�O�ȵ�>��v��d�@?B"����4�|�uӏk���6�b�hw�$[@�y�}�g7M}v�,V�����tQNd��?�!�ct5�w'��ZX4�4On�45��ka���@�Z�#γü�á�~���Ey4҅a,Zn�xQ�6.WA��?��L�
�d�A$Ғhv�� �uO�3y��9���L����_��Ĳ��F����=��ҧg&-�03����K�ӎ��| +Jq)ۨ��
X�u����Ϟu�hV]���ă������1\�Wl��@�!v�)m���B�J) "vMu#Xq?����l�fFZT�;����)B�"�����)}$i!�!Ao �����7�l�R;�k6[ݠy�Y�8��VEV^z��i�����7�U�@L�ټ�� W��.p�:���p���J��K����]|�P
~��N;(x `�1�ۊ������6b�;;��S�Mr���N�p}b�%N	�M��	��	�&��b���78��n0��=�;i��"u.�����e� '�[lR�D�R�a�F�zr��9p�����ד��U?K����>��v�:,���B���{b@��m��,�?Z�\Sߑ52C���� �ʼAc�8�F8i{|�X�$�U��d�*Rx�\�cY�z˅�ADozcǼ~;{"j��Ʌ\�8s�����7�K_3�m�q�b ��syXOl��
��!t����`�����#ܚ�/:�~s�^�����6�������wM}�W���+�L�_ฟ�DK��I�ڝ�2�ǃ�nb�2��P�����嘆'�_8�~���*�G͆�FYȸr��Z���p׳ċ����٭��C�8�?�2D>ڷ��]i��V7�������U`*�Ɖ�b=�->X<c�ւ�ر����p%���ʷ�kPW��\���1v$)���wj���G�����yu��ـ\BЕS�(UM����b�Xzz�7Ooiؽ��!$_�n��@.�"�X�\x8|P�:^$H�Z�����w��� �;���
���\���R%CZ�`X��-�~��{eu1�F}�H/1��z&%G���uh�����b,ZF%�`�Ob<E�/�e=�J�����������Nͫ�;߂��ƞ��+�߃sUԽ��K��1e�v�����"A��D��L	���(�j*P�T���m��d��P�}r�YFY�#D��~\��)I�tFU��slF#�`��m�h�Hx�^�(ke_�"��g��o�WVĽ^.��0�"9��7� �-�H�Y���$�*â���{.(�M6��gv��2t_�3?'����DG@��ڸ�j���Ȕ�m���S�y�Y�O�շ1�D�ٸ�A\m�>�K=�� �/s�r�����/��j$ow��:���0��-
�,6�&I�+ �-ߦ��уԮ�? m
~�F'��� ��i�Di���Ĭk~�{�7��O��/� _��-��;��z)�fu�	����H;�9,��	�{����Y��.�����! +&�f#ؕ�����9�Z~�����2Hfd��_��L瞂�
k߀��(-�5��B����]ٗ^������$��n.���W����H�<�������?3/k?`	h�L�����Pey]�UN���N� ��vGO�c�p{��@^\gȻ���&�oU9ʮH>NIj���`"����j��΄��	kňj��ͲǼ�S��$� ��q���*T��oŶ�ZT�@e����S�蔄�cPh����vnET���J����9���VX�M��[�J/:�ՠ�J�w���!=���#*Z����ץ�.];Olf�7�!�l-�pC� Ġ\��C$���m��g�c���c�7K'ֺ��R=F)�PN����:}���O�,a�TvW�UN~�%�F�����{�p��:�My$�FI)f��p��w�-$!����ɧ}��̊�à���(���E�AF���N�ICc�3|��"-;4fC�G�a���s$�㺳�s3�|ͯxݶ�u[�A��܏���sւ��z�'��c�Ľ�]�d"�m�.�IRS��]����C���������^�.Wն�2)7�yp�L_c��A��_��ԇ���G��PB�?��پ�#��s�9�^���[͇U�6~�m�R'B	hJ|~0I��
{� 5�k�h���"��C�#拧'
>i~L�
��z�>ilM�?��+���I���h?�!���7S����R�6�'nK>4�IF/I�gݹfl%`:�f�T<�W��.�q�::r��"ϛ����PU~���P�W����9��3Ő���f7\U}��h&�x�S����N����v
�y��;�g^۠�,yl��`���ʸv�dK�s;�h���������K�Z�#_�=���I��|Ƅ�N�1�|uC�L�5��ҀH�@5"F�H��DZ�{���9��h��,V,�}]E�y:E��������7�y�'�WB������OZ2���˲3R��B�/o��W��|jǝ6�1��<Y5��.����m���P5Xt�����p/�{�d��TWs~[c3�I�"�lUM�����Y�B�99� �'�[������V:�q�`�\���08�A��Lr1 ���R��{���ueTٮd��a��w�Q�{�<�a�0�zq6�R���ն�=��֊��PM+,��&QE)A��L���][l7g^�4�O�qC�ダ���*�ߥ�������n�V��A���Ő��ެ/�5D|a�_����L��8�m��$�x�d;�yh�]W�t��r�<A;��ߺ�ʧ"M����p��&W�݊����_
 ���G����a2�f(��-�2�z��t�f�.�_���r�4p��u4�/$Fo`z�S�U@��B���U�&ig�y4 P�n�_�u�Qc�W=n/9�h;�6��Ah��X1Ga��M��]�����^�)��kWH�Rl23YI�]��_�)�q�A�-�3��n4W�	O����z'}ї���FV@�]�F��1�Ms+ �<�����y���E.�&s�{�b4���p����x�����n��ǰ��A���5��oY�@�O�/-[vP�tҧZEt~�-F�3�Yz���@����_݊֩���Nt8rK���s-92)j��.�������%���<4����j)7B�k�\w�o�y)EQ�S��o/b�4����fYT��k��E:�IY58\�����|Jn����`M�G�������2�(Mb�ț�G|���F0�ϳX)u��_���
��;�;:�oN��|N�R�6K����w�ܤ���=V ��s"#S���hm?�~�B�c���s-�M
�0X�A	Y�F�#�6�I�T^s~��N���$�}� ��e�Q�%
�߈���}
���0&]l��_��o�ѯ��1�* �1b�X��u%ō���90���?Rwf#)��S%ʔFbڡ'�Fm~�==fb�0��PMᯡ�'㷹��H��F�IE�탓|�fw�[�>X�[ۼK&��`�
Y������۵y���
SMq��v��eo]��=qPw�{��Ğ<>.��/
Rf�v��vms�����*�%ƥF|el0\_�X+��-��Z����:꥝�˸�E���f˾@�7�%ˬ������h
F�U�D��\��^����l�`Q�l���%u���lAۦ��F����}�>��~�;KL8������ oto�*}��-���@��A�vm��m���}玏���w���n�K��)	x/Pëg�u�q������hB�����b��w��*y�\�ٟ��)(3!չfSƄ�u:�j"�� h�?��W(x�|uz���w����C'�)B�``oݺWc��X���߳��<���������P�
���=��/_~���F�]�[�CiV[j/��u\�{��3X�bd��.cP�R3bM��V��K�6�l&�>W.�a���wj�1�ֲ�����LP���f�vt��{(���aHr(_��Z,�9'E؝j̀��і~k��t�+�89��*Z֙~� ��͌@��Xo0��E��X_�������D'ڼ9��c�
C���ˮ��M�ޫr� �C'y�M�1����i������f�	�����7&0��{p3�L�)5a�wu�g����3H	�!��?gҘ(�q`�R�ɇ�5�27|���)Z��P�bp�&4'�V����C�x�/�5��lX��gS�`W���Lz��
6��bQ �4�z�T�����@,��TLg����[�z�PD��%D�%f����ڵ瘀n0\+g��<c�l�������%�7�~N��A(351d���.���)Ӂl��DaA�/����Oy�2��1ƾ,i��2*�s�W.KW;%3x���0ơҽ���A�%�O���TdG6Xs��X�H�,,���ڂh���v+�!��l��e&�%X��~�_��� ������>�5���om����n�%4Ja�P���R##d�6�jG�"*�$��q��?�~F�a�=��wB��X����GK�(������j{��e+�:��xV$��i��R_���w�]2 ;�d����;d���\���[�]�u#.�m����>��ʇ�I�PQ���5{�[T���=i^�KٕP��W*@c�:���mU]6�}�ۮc�i!�W!��lB��C�3=������ǒ��O%�����m�vL�ؑlWG����7S��^����3����)|�Yh9�c��$���[�&P-�u;ݺ�7�R.��E9�@N�� ��L̃3ϧKU�:�����3���N�a5�'�"(�e����OL�����H:>Ó~��[[��f�Uٷ��7��H�Ѐ�G�<���▙�Q6u����p��2�'u8��1�;�����f��e;��p٧$7�hv(ӈ�X��^1��?��:-,��"*U���Y�u�ܐ���fm�Et���}@�T�U	��|*~Y�A$,s����lGf��t�j�u�~��\I���Kt��-En�:�'��\�����c����m��J��ã���wM�u>�]�2(J���䜷��4)�u?���EZW3�]���W������_t���eQT����������}���c��ټ�uؾ×w?��#��j��;<\��({����l|]�����/��a�*w�^�ႇW`�H{�1�4_��0 b	�?V���I��#O�u���}��F7��^ui�����
8�T������hIy��Ke�mQt�_/P1���Q�;���j���K����}�n��X cCㄮ;�(��)D��cSr���%r�)�	S��S*Q�mMd<�����׹q8���q�r�6xx�]��z�A�����7���8
Z�������[k(��_��W�k~b�f��+�,>�2�hWU��_h������E'u���Ht��u�2����7n����y�Hf����Hbݶ_#�F0�o~�}��i'���~`Ct@[�Y<R}���o��u�����2��	o��䩔���+�qjޮ���X��๶9CjLk�3v$��L�s���fWYy��<M�oT��n�I�6V���m�nş�	qMvS(��g{.P�/��Q���?��#�%zN�K�����!y=K��q>��1�<���}:}QR��X����ѷ�����I`b�_�"h�"MW�JX�8#fd&�o[�M'L�bR>��EQr��w�B�,��r3ʁ��ugv��^�)��:�b|ڗ�Z��'�@�1t#;aF���ê`^��P�D�����8�l�2�]HqWa�ňQ��h*�� Wzm<��<yd�
���S9XKɕ^P � ������C�Q�����`4[0 e�o�hj�n9R������v�Q�"���8��}�auT=;wd�_@GM~��W�3���^����<�}G�%�מ��YO;V)Nj� �����AqPڥ��^�%��9�3.)3`MH�������A�r_(Ťy��-c����������K��bN��� ��� �Ή�XG����g�垉��=IJ�:�D��r�� #���1����<<�������2 B��_D�9y��+x��CG�9���X���͝ɲ�<���_���ۻ�C>sb�P�9�bp��j�'f��Q����Ic^�z�����{0��Χ8�fU��҄7ߧُ^.�~p��\=�~�3�O)t|$��FMDfV�!yn�M_��P��C�'���w�x���u�k����(ll:�@^o�z���O��6Ul���)�g��W׺d��h@\�"�@��@d�{F�\�~�h�z�`��(8����@n�~�Q���M����G�q�\�JBr���C���~*�?+�� �uW��g~p�&�sh��_Z,�`������K�W�h��C�՜�|��;��ěg܁+��jQEU��r�Y������^j�<>�2���݈��~h
I�V&� "SRE�g�%��Gm���a���Q~�0���+�!�����K� y艡�$�YG3�P�{��>tdGSC�p�;)7�;iGE������5{50�@��7��hG�_����{���!������1W��w���>�|н�&RWJd	eJM���d�?��K T9'Ņ���-�O�*x� <�-ҽ�+"��s�A.q{��r�{M�-P�	�O�y0�I�u���i�=IL�}v򢎲���	���Ɨ/�P�!�@!�?[�M㹙l#}>�`U�~�$�Lqw�G�IS��] �Spg)���A�c۴��p�@$xB�����ht1U��:@�����#�*����g��y���k�DB�+�l�kx
C�T>cqܰ�Sd��:�eB�v�i���Ƙ���O�ȟM����3��ڷ�!���J�q-&[�[��Г9��TE���i��* ���D�{T���ն#�ҕ[�@<���n�*�8��s�m�����B�2�pD�S��C�lf��a9�,�P}���C�0(E��:��ˌ���C���5��Fe����&�_z�R�e#�%�I�ք*�v�+$�S�7e��ۘgs�[lvsD�i\��6���{OO���5�\!@�Q�T-��<�7-*��n�<<���Ud�g�����)̀�V�,�P��|{>�I�f)�(��ϟK;������B��<}�1<�9���D<|�0�ؔ�'�&�1��0^(��?��.Q3��˩ӂx��=zh�2���4?&��aL��P�?�PQ��o��`�l�L���D�A �[�=D ,K�,��Ds���>@�ޣ�`R�����8Ƚ���t�=;����\�R 	�"�F���EA����<�zLY��G!#a\��
O���j�=�Ӻ~���k��~�ШΘ[a���z�OU-�jY�;${y�ѥ��1--��'_��X2)>9),�k�%�f��毷����]X�𱤫\��y�x!z��l��
��b&�y�e���L8�l�Z4f���3�D�M� �E�҉��Y(�\"ͳOz��#��ۄxԻ�����Ӵ��C���,M���<UX5�%O�ڈ�lo��UU��%
T���7��������_�y�yPZ��$����o&�WvN�%�Q/�`��O
�����U����x�S}0�so�&8 n�R؛G��mz�oOSyND�7�|�a�4ko��`�����)R�ǰIˑH3=�p����R�����ת�xmm��� -Y����� P��>`�0q��0ڒ��xo;�V���զ;�i'Pg����ÈG���[1Fw��b������%���/��!O�q�*�o���u�
��+�$�F��tH�گ 1��X������?_T�'��`eR(�ebSq�g�Z�nF�y%邾�����C&x���kU�����ܣHM���9B���i��*.�*K��s�dЖ�\q�ڍL��W�����xa�w����L�����̯��R����N��������5��s�I�X!t��fU��2@�Cm��sN�џ��X��x�*KO�3� ��Vi9N��� X��BOa!>j|c"�}&��if����5b�C6��j�ɑ���=%q1#6�˲�Ȉ�S2M5��H��8���	��?�AD���u���'�,t�&��`Y����}�:���R �W������q�<�eeG���R3�����l:���$��$ٟJ0`'�����	&�0=�ⳋ4{�@�d����&�u���.�-�/Gz��K#.�rh��",��'��Roa��?�0`+x�@�w��&��r����;D�h7�Ę�����{�I�����k��Vb����%�ט[M��7$�k7\�����A�	h ��D��F��.b�#�gu@��Gx�<PC{>uxK\�-ፎ�*�k���;އ���]+0��^��8��,�`;X�qi\��/�Q�̶
aRa�X����㍆47�Ym*��H�KW,O�zY��4�˜�H��^g���A��<��)�����J*�Vs�}:t�т὘��e���L1I�D�1y>ܤGK�V���ϩ�2�OCP��2��y��h4�1��J	qīCf��D�Fv���`�a��	pX�} �U�q!�����LZB"�$�f��?��<�8k-9���S��9GҪ�Ԝ7̠��C��p��.���6Г������=�>�p��RQ��7�g�e�:?���|"w2��h&m<3`z�q���:�B��(��c|�w�Qu~R���F�7�L�[6�C�`���<~�0f�W�#h�iy��%<2�9��L-6�u��F�pa�h����M�] ֪������i��T� �z�� ���B�coV��Z���[U�k\ub��/�HrA�ӡ){QSt��ZfP<����T��1�{�����`�/5K�<�G��"�]����,��s�c8�'�\N�pRu-�x�6�����Cc�O(�e��/ŏ8��ZD��V_ߑUD�2��E���".���$N�A�t�j�)Y �_���՝/�&�+����S	٢����g�TE`Hv's�w�c��@���K.� �M�9�Z�T	�(��g�Re������!����6
�?+'g\�d�G�par�y��T�Uz���ɚ\�T��l�Hh�h�}0�쥝��ěol��+�v}�-��rz��6={顗ƈ�+���R���!����+��}u"+�Z4�<+SV���ό��7��eI��߮hg5{ϞJ���	ZҰ�跪Ȥ�� �ݡ7����;�-��?+jɌ;�������	'\8�Y�����5%��7o�.t�~2Mp�a��mB������nd
�F����c		\|]�y�jn��&}(�6�~���O�9�H ,����5V	b/q����$��9Č'���(9�E-�;3�+n¢J4��2�q[���&�#�YˌS�/_*��Y�aø�s�����i�[rF5�[[9L����@<�y��VZ6Z(P�M|)��L��*g7�2�2�WD��̐���8����Y���#����+��M.|��+�Ay���;����X�faE�o'^=�S��(�$�Z����B���>Ξ9��v����Ih����f�w�rS�3��[�2��` UUǢ>��GB\�m�zx����L�7l@f9��"M��_=�
hv�1Lr[��6  xt���7C��^݈�\b� E�Aj�4��ʨsy����.�S�z�8��oZ��Q����������#O����a}��~�o!����׺5$��Gb�K�����hk!���]�������� I���:��H�W�B��K^����>�eO����?�DKI��y�?I�m��x��� g�@'}I�	l����闁�H{�9�[^�<��V�5�c�C�T�����5/�Xi�3c�WU>�~��u�����[�����IE��I73��ZS�G�w/�+�i�y��u�p�"�E�N56�2��#�}�4 ��-�J��Ɵ~	{;��^>��X�?@��!_���|��@��B4�w�-�'�cm���B���+��HI��wD5:�.��
���7I�!Ϊ!N�Xԫ3�t��Xf�͖}�d��Xz��KHX��|Oˬ�� ��D	AHz������t?θ�ߣ�>h�\��A��<a'C(<A:ݏ����'	��	aj=���Q�N�~y�|`��'�-ޢ	��5�^���6�@���&U�ϕ]��JG�O<ѶwV��L�$8�����Q�ڂ������`g� '}	����̃krI}yH���i�Q�C�g\��27؏;ռ,�{oY �P/�������$���Q��1O�M*�*fi��7I_���Š�1(� g���-�!�;��ǻ7K���~��6�������|�c����m��B�� '
�~n��X��O����w��H��;�9 �'+�=>�y�+�'�d��0��`\�U�3���>v��#�õ�|��3f&��~��	�6��t����(����rT]Y����Q���O�ʁ1p�Z,�r8��t?ٸ��*A�D�G��/���S��!N��W��y����Z�����|̝���,i�x��W�a��h2��4=��߿?��ś���`0!����]�9;!�-���iC�J,M�MY�}����a�gk20C�������:���: �RvFH��:��eD�*�|��N�zV�dpP�I�,(�P�xKs�Sf%y�?I��-0=�"�!��4U�=u��w闥�ܣ��/���:;��	�Q�� ƫ!���U�V���e�Ɵ
��O󉦸��:��j�AS/(-���rJd�ui�c��>��Ԣ�IK�4;��	�;��j�zu�y���Nh���<�^��s�>] �������Yޞ6��V��D,{�$�"5
4@�~���p-�z(2�G�A�6�E^7re#
���)�ِ�6̹K1�O-�Hƫ94橇�����3{Z�@��޹@{⌵��]��.�2.��p>aҐ����aO��;��~�������̨6�~L��^2�*	�I��c DB#��Nb��^��(�j�\n�5Э�,�0n�S�qw����y5dǸ�/��GP'�W�&r��k��Լ�ϪE`/Aq�0 �_�'��c�Gu��:����'��%����r������8�u�br@���ׄ��@|/k��ƗRs�����)�;N!ۃ�x<��Q/_[�7��FB�@`�!W4������Mdm�Z���5���į��Җ��7�7Y(�99�(�= ҇���)3}�����y�vˑ��:��mN�觎����QT4��N;0�p�K�e�8-�m�Wf$�"�
�Z�K]E��/)Q������鰢I�_������P�W6��*%G�����Z0�������C��~����I��X��x3��tC���^�QCN�Eu^�_q���6�{��U"�2mxW-��og��p��750������ux	����O������Lwqeh�	��NT(����|���Y%��!��1&Ǫ����rp�t��m�=��/:&�\QXvg�AC�/��;����|��':�4�#�IT�i�J���w�0���f�N2>_��h1v�]�J¶�n�9M���{+	�[�#I/��c��X��a�4��$���c� [-�N�*������)B�Vf��Wn��aAg����֩O5. Eq��J.5��O����,'8�f��A)'ZX��U�	��
uƁX�F}�>�]��R�s��2w�7`�5�������/��>�ͣm4G7N	��$��x����w�`�e-��ܮ��<V2>��8]���f�vx���p��x��'ֶ�x�Ś�8���Q�9��w���i`>��iqH�/.���p8[�jVE1"�L����.�
U�(�O�B��u�����8��=�2][gb�����Xژ!?W�^jv~̰�;v�ŏ^�z9�''��-�sb2�[�;�VT��C�Ҙ���Bƚ��yq�MXU�u�����|(���ok�������y}b�Uv�׋�r�%�v�(_��eη�4�Ӷ��C��^4𕓬7\�D���r<r�,�p��Y<&��A�VS��V���]ay��wV�k۠��SI�?�l��3��	�5^��Z"����U^%��k4�/���q����q �}a}���%�ւ�߇�E�����ռ��c��v�S�M��|ׯ���9�`z�$2ѱs��|JJ�@0���K�H8�����|��#����x�OGó߮�G���4I���{��K�gX�?��~�1�_NmA��2�d�����c<�,-�x�7Qŀh/�}����u�A�y���)�K(���U0�V�#g�۪�ͧ�"�4�Gٯ`�����T��$+;��Z`S�Pw���		ko����Ys�<L��%X��ڗ� ����H�8ןA�
�/-���6�����oD@n�������7d�Lْ�ZJ��g�8� 6o%��ퟫ��fDq@2�KD�u�Q�]!0Fqz��x�Y �͓��f��I<|lw������_=��r���d��X�%�ق�r�Y�T�"<!�2���4�Q���������5�6�?�$�z�Ď\�ٮ, ����=������ ��T��u���5Ӥ���8`�fz���|�n���������7뀦��T�Ƥ��.�
��xsi���e���XB,�{R�t��5�o[���t�%h������I�cf��Fw���J��۲1P)�>�Y�X���Y�+� �.��m8��.��k$ߵ�����}�L�)�\��}{�����Qs�����J�(���I��׼��-��Пv�Ҫ��vPP8��Bv�`�Q��j^�!9P>B�6h�B )���%6gI��Ff8n����	�Ň�rii�����s���C�}�{��m\���K��+m��.�SB��L�ڵ�[��D����n��X6l���9��nO'����J�q1��\��F��CIy|~����)���4f��*衂�[��2��r�~u�|������;�ujy����Ǵ읕���/XDD����;U�+��_��n$�S���vv���T�����X"�O��鈬o�74�E_�V3����x66D�`���N�*��e�J���+1³7�dFe�O�K���Z��H��/�Ff��6��"�
j��\�*�bI �l>���o&����w��L�b��6�z>9�����00�#^�Kdґ��n_�:�ec�����ʲ��!�T���w��Q���]R��b����e?;�m�I(�������H��)�ikU�\�<)����t6x��l^T����0�u� 2B�G�_\�u�w	E�v�FD&�"�
Ƚ�H�V~�:�h<|�7���Bg�}S�L%fe��ܤ�L�p�_:�=#��J�x�&����ZL�ߌ'���B����W� E� 3*�ﭥz�M֛XQq� D
�7�r��0E�q����UJ����Z��<;OG!F��cVY��B&��f�n,N�B�ϣ��׳.��;����澸�7Y��v;�������O
M�L�^��)[e��1$����1�ra�G�i��*�])��Ns�2���e9:���C\�����ԅ=�+G2"w9r��F yUQ����p������?8�O�Hi؞�z*�_�b��&7���R~4�9O
(�_�� �L�!�6*�h�����h�g����?�ڶ J]�f����g�LO��v��{Si��@��OU����60DI�~H��\���I�u��^c�.�XM�L�$�qm��5w|�[m�6ak׸�R�}1����_Q{��������͌��2[y��-��J���&��f%[��b�N��7��R�N&I�.xH.E5� �����~�E�c�"*�ϩ����udcB�%B�U���Z�?�Z��5�Tj��4Ns8퉹��U�m(Qy�5,:��]��\lp���p�,gC0�amo�y��[ϰq�p��
/)g+􇙔��"�J֪%�gs�K��fKU�"���K�}�#�I������u�D]J��V�e���?�D�(�W9M�Q���Jq݄��vי	������\;��3>�Ə�
�w���U�G(��u���C����ׇ�V�r��(�e������0�3�B��AeU�|�g
E'��OL��_��F���=i\�ĝ$�[�hC�u�hM��KY�ڕui����J�Tie���V{�
�u)Bu%B�"�6~�U�:��r�|���}f��y�����m��Kk
�գ��B�~۾Գ!�fdk��4=��v"����9{�+��by�F}�l��x���C��.(��ܸ�
O�1ݚ������w�g�`�?+��Ƅ�����>�����bUb��!� ���QJ���[�q�Kb��[u��Vp#c�;z������+���W�����ͬ�S��_�±�"M�C��o������*0�sw� ���j�v�-����>yMg�n$��|⃸ti��S*i\��/���`��ڵ�=�����g�d1��]�˝��xU��&�MG��|�d�>�+}�ǃ���b�ya��̴5��%�˟�FR�n;E�#�v�3}��ݚJ��Lc5?��V�@�xP`����-<� �`WQ�x�S��xw�M��sA�FV��&�x;C �*�*�V׳9���p/\)��ƨ�)��#;���q�x��v��z�K�u�8�����I�u�׌����d$����z}�i��+{�ǁ��R{E~�F�5�@,�N4��i_�ǫ�о"�u|WR�dM�`�I���`$)�B�Ճ��t�\�^p�3y"+H�9τ��4�n�E���C������Upm�ѠQ��U����ifru$-���f�Y9o�g�,OKa��`����-��L[i�c���B�=�a����3�{6� ��p����+�r??,��=wh�z�c���L�Gf+u������A����zKP�C���A��Q��!��x��f�qX�5K�<���/o�0���85#�ԝ� �����S۞����8ɚ��u�-q��1h1Y����+$�c���V����^�d�E��Ñ�.�PI�!q�gԥ^����'�V'���#m*��NWC^��[��!��#F̙�;�w�$��mf@>�����y(���H�Q�U��*���Y�*�YԮ'L�t_q�yЯ^�,�Ɖ(��/�F���P��Q��3�m�䮹�o�}K

��*�uQ��2���+L��WN�A����0e���1�٬Z��"�cZ�n
J��g�R
�����F��B�����o�����\�XM��α�e�X;/��c��@���O8�ic��P���(�B��+;�ʗ�]7�T�u@*"oG��������s�\R^���̲-�8.��-L�GeT���R
�ˋ9Vs������Ŀ���:�d!�kJ�u��q�E0���.[�Y/��^/}��󮘾�R�ܓ��P�V�~u�?ö4��5A*���Ɍ�����<��Uhj�Y�;���*���)�c�X��1�U�����Z1g7�p��#�1��U:�C%�N��5�(�cȵ��񦰈?�ӭ�w�����������䵔.��p�h<��"(/u�(}��
G�g��T�[�I��H_��7�A��WlK���O��,*Vh_�Pih3}�7_�LM�t�hZĽo��)�-gI`��?O��W�Xf������^V���B����S��j�y,<5}�W ����'�Z��+�ψ@]KK��Ci�ۑZњM��/��*L�r�>���M S3�G����	����`d
��P�O�$��L� ���4�Ó�3�I@�.Α-S�2���i艶ͥ���F�T^Y�MtOL�+T#~�	�W�����!�P�;_�7��~���]��X���5p�"�>"��<�+����i �L_ظ�Bݬ2�v��ٳ�[�ޅ$�-��̬7���5X�~$�s�ʓ�C�����y���A�Fn�e��2����,JI6���.�
�t�Ø_�����0�5Zd��θ�����`����<�X�<�
PN�i�p_?�WK��~x��?�qO��7�P� �������oV��'��=�Ӯ��_����gDY��%�|��#��c� :sv�5���0�e7��F�%�|��kZ�)ʘ\�j}I;z��RvM� �eQi9�==�Ǌ�Zym�ˊ��g1gq�y@�3��c��t#�Ky� ��oٗ=0Mq�w�MY���ݩ��L9�"D�m�>3����[�~�8�,�M���^��Be=�	��'�~�8��F�D����}U��G�_�0>�(CJ�j�{�Ǯ��$��H�_)�V|����yo�,���ԩ�0fT��`J��w�	w�¹��u� ]:Q�뙏�ޛ�0�w��X�����|��k��	��%m�@��)�W��rnU�ӷ��¸��m��]���ev�8/��2��«ǰ����S�pK�
�q����f��>����%H!-G!�����/>��ok�M�xt�՝_�~K$j=(�PK   ,��X�u�Q�"  &  /   images/87392e8d-b818-4203-815b-f0983b827fd2.png�zwXS۶/ҋ��RC�H�@���DJ� !�^BQ�I�*E��H�� E @�)
��}������{�{����oe�5�o�9�o�9֘I��(ə����(u�5Lp�-��HJ��d��r�]ȼ��|��(��kxY97���v�K?K���H���L��»:UP^PG�� s�{(��t p'%�������:���36�8#AN@e�"J� 	�PHw_y�����+�(���T�j X��=}` YqaG111�,H�A�Y�H�I���K��KK��KHˋK�<���|���M4��9�I	����%/*(()���"*�D�$D%$�qa� ?(J�×�/0_G����p�u���S�T�w�O��2��L��ET\DL�/(�o�W-�ű�_#QP�:9�����q��%'GQ�;	����a���z�z�y��z�7��n�wK���g[�ȿѾ~�~�3��5��z��8�4pfrWdɫ{"�|`��8����
�����Q���C�A���H�	1���)������W23���+���(�����?�����&�j�����K^���i�N^+b���	IyiYyi��br�bb���{:����K����ؿ@q�8A���G�������s����D�<\���'G���n`���먫�x:��qZ0�C����+���u<|���0% N"�;�KJ�88�ʈ��de���` a&#,�9�9��KJ���_����*�������7�4u�_�J.h҆��y���tMa�޹���<��Q��9��������+�����|=���>05���8��& !)"�ׇ:�=�$ust�z��p�U(�sG�?=�w�E�-a�%�e�?�%`���)�S�KЃk����8>�h�AP9����>��u���e�@��Rf�v���qe�N��iƎ�7y[$W�>�p������It��F���MX��\!ȧ��7B=��#%p,�c�Fs����'
1���~f���NZ&��H�s�� �	u0O���R��`���	L�پ3�Y��z���o@��tr&31�m�Ĺ�oAX�V�0(TμtL?6)����oM0)����F����G�1�M�g�0ؚ�گ/��,2���؎*���<tQ�܈�vC3�]_ָ��Wn<ٙVJ�ҥ������a||�}_]��SV�Y
�	ܥ���ʿ- @�{"r�~3�N��,��m��m%ry,�|:��V��))G��w|���e#,��xM�ᯠ�בu�T�8K��-!'ߢ>g�
��A	ԡg��b�0��l�.ވ�"���:�8�m('���x{����qQ�~��j;��2�!no��CU�O�	<m�~�)\�U���ƾ�w��C�� �F���B.��ڽ5.��߼{]p|��W���m�`�H�������;jfv��4�[�������T�$g(��OX^�4QG'��LK�bP�
�g�Q�s�
����B�][�~{LEv��W���t�y�V,�)�8��1M]��PM7�y������+#�ݴƙn��=�&['1��-r����C�G��ޫq��ö������c�g�aq8�k�}��
���F%�`{ycF�8D�ԧ	FR�����-�3]ي9�ׇ���W��j2�컑�ґ�����u���&&F�-:M��N����wB"'�w}Osp*(���$K����?F���<�c&NӢj���n%@��w�b��ڎ�Rj`y�L����Z<�L4��,���֐��Ţmy�V?
N܀�&Q�����Xqj��+�:�r+��`A0.@��1�w�"��)���X��7	�v<f���S�h��i�V��J=}�����d�uin8}�掳��췹+ݨ�!^�N��4�����Y��&E}I��˸Rr��wӣt��1�����72�����ҡ,����_)H�$V܌Npɧ�'�tw�a}C�:>`_��j�?0���(�#�bzr!�X��F�P��bD�|�ݣ��MT�r�Oњ������ߴ�k�o"]!��A�tE�ʱ���~��i�8|g5ܑ�D$ �trZ'؂=����3��O�����2��-vn�r���^׿ҳ����	������B�R�!y��o)P=TQ�c����*M��N�<k��EMDT���}��~S�( �Kms��j�2����8��F,�G,V���j�Хld���H1�+d���`8o��������:�)K
�a^[�XT۶uO��D��1�v����*��7��Fg�{��k��"Z�4��
p{�D^6�t>;U���3������r�%r�UU)s���J[YY]���
�&�\��T?gY� p>������64ܶxs��p̰�)��V�L#�=gzbb"*g.@k*�uq!�]��B� �k��ZKwD.V��A�ì�CzY�sVi�l�8ã��4<L�w?,E�Z|�����z��4��.1G$Ǒ{Ě�M��b����B�I��4��?n�5�+���(v����al��I�^�����4�Hr\~��.9���3�#]���/.r���^i����5d�/r{Tbd�� C�n����KǍ�U��9kC�z��Ç�^}
�l'���I�[��q�ڂ��^0?1I����hͿ�,��	�m�6-�����w��W{�R���1C�dtO틥��UUO>���.�|�'XP��5�}�&?AA�FB11����%+[�tla�������S?MZs�}���R����-�i��$S����4ת��P (����-�c�A}�\�Y��ݷ;�CZZZ��\I�!�詼#��%����=;吝�%��Y��S�l�SVèF��e�>������u��ZJ�$g�;��Ԍ�<��X�ԷDv�yWd����(&�9���i����}8�!|�̦p��Y���r�A(��:��d0� ����"��Rq+u\W*��=NE6A����|��X�sm����r���M%3�yx5�h�u���������vYn����T<���|�(�kb�7P?�`}�C�ϳ���®��_|��ќ��Ei���R.C��CY+tܐ����V�+Vֶ���/<�9��T��񽙏�E��˳XlD� ^S�F�~6ӽ&�d֛����z��u�>C��a;�ikR��� ^q�CNF0�L���V���/��-PF [ ����9N�G��M_)� ׾h���A����[*���u��f�I����s��{��^�J�vU��U���Ѫ3g�`y�b�#`f��a����P�Q������.���HH,ԅX෼�|�u�\�Is+��؞�E����4��\��]A��r9z:7 OW�Tz��Vx��Y5�ύ�f�.����P�b���1���P��M��qZ[�\����5�gkEZ���[�A4L�������h$���$�IA"��;��B7�Z���<��������ý`�F8[�����֡*��>��l"n*�T4�3��\�(V��L��ԇG�~�/9���T��{�a,e��,��<7r�s�ҟ��5PGj`$g��3\=#y�6B����C�(����x��Ҭ���X���*P.����#n( ��M\�zL������L���qcZ,3����7B����f�ucXd��)���
��S@�}�*1/���'�<"�W��08]��B�4>~i0I��*�h�Z�ҧ�+wcΖb$��j7I��.���p&ବ]�`��w��и{�@G9�[����Ac
ڌ�BdҐ��17����mk�+�I|�iB��	��ڰ��K�[�)覘x
��]U���^0r�ׂ"j�)A�����E��^�|b����e�8�wf���UL<��VR��Z*�[mCS�������{%��9�Hqڇ�D�es�l�e�WD�[ʘ�6i%��.�"�B[h}i+�u�P~��/��(:d��������ϞZ�7�}[c��>f�΍��6�!"z��y��+��u��9���V�p��;�����y����\	����מ!`����B;����_���Qi�t#y$���I�rަ�4%�kt���:���')6���h�a��*ǽ�>i�������j��:od��*�q�D���
@XM>&v��0�!�)��%��׾�wAޮ�̎���**����hkB�Ѧ)�x��/9e..�,D����~"3;<�d�O������F?W�8�����'T�(t0L3��[~Ov2*JMIӸ�̈́�>cy��bj�Iy**�`�Us[Y�|��ME��Ô_��B�<
���c��7XB�㊨x��$n��Z�㖧Hv��",ܻ��˿��0�#f����l�k��(L�Y�W�ѫ��cޮ���\�q����T��VONŭ�6�T*������w�֭}Y���:98
=�!~h�I �� }9v�)�����̩��c3Fހ���߳�'��h��b���9�y���Y�V	+0eO�!�y�»����l�<氌����f��>VJB�-��A�V`�h.s�r�f�|{�u��r4[�+�#�şͣ���zVI8�6?��� �U�[����uj������G,R�'�vp0ܷ"s<_����W�͜��B�;#�a�aw��k2Ebg�ƻ/$�����{]�<|��c����|a�N`"�\�]��O�\�2#�o��/²���$�����x�30�#lB\kw�W�O�LG�~�I?��g>��k���7����jM�ȩ���Q_�.d�r�x��������5=�vY�%�����]�Qשd3N]0c���` �s��C2����/U� F�)��]Tf�~��b4���ȱ����pȒ���_�;c4��xB��sB�oL�Z��*o�C��I�.3g��2�e���"�{�9/�� V��&:�M$3�[���"�G�+����Q�n^��Lk��uܞ�:~���h˯��J�d�יɉ���[g��ׇ8�mT�%�I�hE������|�N�J8�#�Scc/��'��M�Q�=���n����އ�oo�r��#��ϲBO?D���+/�\J�]k�U�7ڔ|ů^H�v��.�W*�H�NY��T�t�һqN�VO+�Gi.nk�Է��V����si�44,]�[߀[oI�y�i���qF��
�%��y.��>��I��̃�2�d��Qt�+tX�7d�7��5=\2��q�;�[�[����m�ǒ�˵�PIV:��YWz����C6�\�f�������U�E\�苋���-�l�Nl�T^�'��ƗD�����#�H���J���,I{���7 ���g����]�rŗE�7���O�;��JKK+8��<ѡq��Z������^6�!m:QKT|�m����s������I5��6Sa)a �R����� �xI��q��8
y� j1���F�.U*�f���\�1��%Fޤ+kk���I!�O��7Q.�����D�Q\�����z��J�2���]9t�3�,mHN�:r�ź!t��'�� 	l��)�RN?Q�׍�s����WS������y�OϾ?�T��)N�S1�M��>;�
�dW�y���C��^���ާ��ΐРWj$�5,�'�2��[(/u��)02� �Il'-�!�j� �7�w!۝�h�۷;���O/Q4���v�"��]U�ƍ��j:N´��6dӶ]�F�F�51t�\�jM�4�����G�3�6(���pB���lf�����U>whӽ\�B����+ܗX��j�3cg� ������֍�)%�K�D�3�Do,��ҋ�x�	��d�I�x���b��|�+�����V~������Ri�j}���Y#B+�,s�9JPH=]㝊����2Y����_'/�Z�HBIH;a�Fj1�Y��T9���'�{����#w��E%޴g<d�� ��w56ʾ�����2�&�<?�ɜ��64���?��~��z<0���}DMfތ?s,L��$�#���;�5Ǿ�W�&6��#M�%Ƙ	Z'�Įn��z����F��BL�����|��$ �\�t��Y9�! \r��� �Wٶޔ����R���!���`��5ns��"��:/���3�O�CE��5q��T�Ѝ�
���T�3��*~��K8Y���	]>��7���X\�l���=غ�3�6`���X8��$.nI��ۤ+7Ӵ��j��Ȳ2��#fD�z��&�����:��ɗM�tK����<��}'/�zq�Q'��_>��_�W��}ͤ�����AP�F���=<����]Fȉ�����T#�#K>�ҥ�W�^���}`�(�1�HK��u��_�*&��O��x5���N3�8l��h�a��FK5���֓��;g��I���MY���B-�䨐�����&�@<x/v
zǑ��C�Pu�z�:�϶�'[#E�n�D?t�W�n���é�"E	�c�0�ց۫t&�k�o3�)L��8�]��z��#|��ߌ��\�3�`C���v���%��E���G�/��ށF�g?'*l_/���z=�"�L���[�S��_�]M�O5xj���W�4'L�\
�|'YՐ2ۂ���Rl'^���{p�6�8z�At2jb��h�|N��+((�2�ۺvQS�デ=�Ͼ7��tŔ�yW��q��%�sk[�Bf-�>Q�=&qif�u�=�����U��:A���]d���m(�RD{��z��g6�9��R]QyWϬQ�U)��p��pÂj3)�d�W�8�}r��N��Ni���(��oM����� K}�M��Y���a$����P}���0q*��� ��|��A���R��=�d�'�������Eo��F�fSe����̹	-�����ɍ̲l�n�RT<2���E��2io�x�6/��?q�f{*}�bU>bD� ������� �G��K�)��6�S�֩�����Ln��z��
M��s��^�&d)]}�L 9�u��S�T
?���ӳ�|.ݳh��$�tr����Ȥ�?�گ��E�=��˝���S|����Ɇ82X%�TƳhlG����	�;�}$N${�ӧP^P��&� 9��c-贠����3Ao����e�g���PEƼP�I�i`Da�����:���a_q1H������xS0���E
	w]�~�O�8��Vu��h�?�i�)���H����_��ԭ�C�+}��H�Ѿ�DXd�`�>��&*�_a��ި[_�؛��iO-ڤ4no�o9����u��f���-�Ǣ[.2O�"3�iA2�򛙯�γ:�)P�4���G�YB�#�8<���?�	��.�n�E�%�i��Xۮ��ҷZ&���v?b�~uI����90���eb�ԛ�ٖ�Ơ�)���t�{�̽�64��w�O�[Af7� ����>&p�8���ڿ<]� ���X���;Y�E�U�'�}F�>��2c�>m+�a��닅�ݡ����1�h�n�w�U�"6~�@�00"d��Df/��p!���V�z�b��x�}C��Bzg���\8�G��ϰ��%�){]*�p�@�4X*��C�˾�t&�?W-�E��Λ�N�OXh9�~8�;{h~�����Y4/��Aa���w��B���9��o{E�H�XЦ��m~��=؆�PjuI�.���u��{RSn����~j}�iAh��u��?c�ēõ������E},���h�Kjfn�g�mKDqO���I��kA�K(wNL�Z	-�R�^��
6���G/a��HG�������ٍ�/E/�^��[3��N�Xb �ڼ�g�tqR�y+���>���X���E�#���1����ӞD�J,x�s�����(S�U�{Hp�����:����M]�E2�����e�[
s׉�F�آ�/����wb��nNW*��u�$Hh�S;O2���dp�����ರ�뤃�����~+�w�����r��FRI�a�8�)��Pr�����[�}k'�3������U�?NX2�Xï�v��'��H{V�VV�Vz>��J�]鶵S��T�zWQ/�&u��I��&]4�xe�rT�53�.�Mh0�� �o*�}�|���d̬0��]h�p`���վ�ܻR!DRU����!b�F�������I[|��D���e�����h��Tч�`q�*�^hP�1T�|�S��H<ق��$u��Zj�l�+����f�ɶX>�Ņ&�~۞청��ZM������ڠ}[���Y%v��_��o/lx�8v;�{Q��cKQi]fA��Y;�IE�ֲL�������j���!�����U���55Ɇ&r4�?�u����L�ro�!H�V����~�G�ʴ����ajjM���C���Y���ީ�K���ׄaaa�$6�k�x�q���R��S_��L=�w��������ӵS�|.��W�ɉI�"[�@l�'|=�VԦ�q��Y�?X�(����Ti���ÃDM�Ɨ�?h��q톸��������C�T:���*�K��Ξ)�?����ښ�|�"�>��el�}rt��Gn�� tQ�eU&e?ol=�2�{sdn���8?���8�^����/QA��W��L{?n���D...?��to����}�/kF�UWW�l��
D�)�%iUn��o�/\.�˭�f)���%!���)� ���۞%������vHa�E_a���3��Y]�|��KM5+��p�r4SZ�Ǝz��r�	�6��Ӱ���,��){5g�r�	��0��w�ј��?�.�M�ύ�Y�1��NҎ�Y�~S�9Ufj���]�gKG�@��>�? PK   ���X��/F��  ��  /   images/906ef243-ce1b-4f5e-9eb4-92ebaa7c38d8.png ;@Ŀ�PNG

   IHDR   �  w   `�3�   	pHYs  �  ��+  �RIDATx��}��U����קd2)$@� �����T\�����b�����E,��P�� ���R$"���H�(� 	I������=��޼d2d&�̲^>a޼y����{�=�{α�o�oc�o����7������a�mlpL�X�h�2{���;��C����vuwT������M_r�G.3#�7���{r����S�ryJ:��l6���^:���4	�V%�;���+����_��W:�݇�xo��<^�̬Y�h͚5�������|�~t�Yg^~�Qx�����n�i�뮻��<����Ţy�G�iQ��8��>��J����EG}����z�U'�x�[c�[�0^xᅶK.��w/���S>t�G���_h~�c��ܹs�������2���$��r��U�VA$�ʕ+m>mg���=����}���a�4I�y�w�%�\�N8�����{  �"���ðx���Xx�]w-�߃/�˟�袋�ݒsߢ���/~����2�K�~�s睷��OAX�z�J�P:cӚ��3[M�eT��aX�:�Y�g��]�����y_Zh>��C�O���3�������y�{i�������ۿ��M��ַF�oB,�H�;�:����x͟����o^�/|�7�cKq�-B�?��>����[n���V�s�=ȶ]�
E�811�T�O�G�kS�=�����p���}��ߵ�#�M�_Yb��GWg�(֞w�9�����O[y�������%�a���i&�7����'���3�8�ܟ��'ߦ�<6;a������΃~~�y�O}����I�_���~�dSG�'�Q�t��~�_�۟�̙���t�9��KO<���7�p�?�V?�p���[�x��)8���8���E���i^s�5�~��o����1ڌc���W_�3>��;������~����W�d�!C��Ü�cvj��5Qlx�4�+Ez׻��'�x��k���eq��%�\�Cڂ�Gi�o��z���;�^���(0p�DI���QVL_��O�����f#�~`���8���{���ݱ�ڊW����5oGDF*���6zF�^W�"zz���6���S��<������k�|���?�����Rɣ�O���F+8��Htp&�f]�7,�~C�al�`�#�J柿��������AJ��S�d��XB��@N������<�0`"��R����@L����4m�1gΜ%�C�b}Bh�H��燿�c�l�6�(�_�hQ�����	��,�q�Y�����6�=���a%�f�����,�u(m��^k4�H��T��(�ʊb
����>�Z����~��G?N�q���o�Ή�MK,���Ot$Ću��j��q?&볟��������r�`y��~��w���[y ,�G����dR�_�@��,�I�:�@8I �bq����s�Y�r�i��}������?!4/��%N�f�)k(\����?8� ��9�y晃|����r�2j�h9a�t�qןq�)4oގ"B�@��⹖-?+�
i70mlݒEM	a$��d�w���ݎ>��c���_/ᏜH�a|�+_9��/���KNwB%��"�5A x�������κ�?�j�h)a<��s����{|���Z��+5�>��w�5�	b#�⍬�t�^���H@H���t��O��s��i3&�����4��$����L^��%K����vۭ5f��0.���?����B���j��ƺ%+b0Z�p��'�e2._���}�s�Y_����Q���_��'�l�$�h�����-3�[JW]}�	7�t��=�V�9E�w$���R�U)Z�`[)ל�j)a\y���$W_}��4	㩧����=�n���;f)ŴYG�)�3QA����}��ٳ��|��ߟ�{k���Yok�!o��④���Θ={6������6��ʛ�c$�����s��丆u��w���~���������`%&���"�E�'�x�Zqݖ��z�#|�p�χ��(�ٸ�b��9�ݬ�a�
�,�ŋ�e��`%o�scJ��\��w��ElOO���'''�Q�eaX��b��R܈^t�A��CصU���|;��ΫV��@<��cq�i�5[FO�����9waÆ�o!=1O7���''X�Cs�8�9s���gvn��V�X�GBo��Römѩ@�K�.ݱeץ�cƌr��`��6E�Y��&n�vp9@<��N��ݴz��Zu��^{mF��zk�D���\�r����n�k4����n���v�A	�ʳ���Y8�r�I�1���3Zu���y���	CɾM��L|D���I�ܻ����fx��&�fs�&+a ����m���B�44�u<I�8u"RxN&�����e����(��0h+�u����M���{����I<ĘDb$��y��f�ey���,:F�Di+G�y��l&�ɇ��,�Z5ZnK&hnِI�~ɢ�� ]C������G�\t8�@��c$��pQS(�b���dA��fc��|f�@�1"[[�4�AFK&�RQyE1��5���
����300H��J̈́*�O �	W�8��H�����?1<����Ds�K���2+-�}�hp����f�ϙ8��3o}c}����\=�붌0���Z�!#�-8�4���A�@8q�v�����^.��.gC���9���r��	�ɐ�$�0 =��,˥B�P�c�%�#�$
�h#��l�ha�p�+��P)�d�-�n���E��b�,�q,�cK/p�;OVrVK��q ���4�<�!�`n!��rU�pŃh'1�To�s&9��$�J����i�ò��G�iG���pY��J%l�ǜ�䵵A0�6���@�=��N�)�O���;;��B��){Z�D��g����9xUIIĕ���ʥ���N�9'��9ژt���D,�)r�J@:�E]
1�F�o ���c�Kϟo��_��;�h�5�6�`D3�T��{"�p�iӧ�?��:�5%�ϻa=�S�d��-�-�1�'@�mSM$.rȾ�����|;��|��fϞ]?��w]s���9q��xԑ�w�GN���;�8ꨣ*,\^p[�nV�8X�/��ne�F��D2�ň�Mx��t�mw�׾��2�����p���W�"	H[s`���[r Z�c���ğjU�=t�O��m7�U�t3��4>�K?vʩ���k�������~�/���}h���{�;��v?&�4+���=������7�y��@���ض#�H�8o:�pL6'W2Z�i���&k�*qpHM�G��_͋��,:v��W�.~����¯��7��v=�����8�?�o��Ƅq�㤎�5�/)�9L�n`?�tJ�D�����f�6)ul@rj�i;�/��8��aۺp�O�-�e�Ϋo�麅�v���+���/���1������ʆa�`�$u4p'�d�Ԣ�-�N�g2�|	��d���c��W	.b�h��~3�h�X��������q��_[�^��/ް�N;�:��!-�Gn�V����c`4ńZr�͇��)�dd������;�v�u?y�G?vƒ���g}�/�4o���Oc�������;bƮ�5�p�U�!�}$���%`�W�a�7w�r�/��r��xξw�}��]��/��?劯~��Oo��дz��L(��BVV�M<�8Fw+���	#����s���=������Ww���;��e��Ѭ*\��u;I8���u����%�`����1��m�}�{�\r޹�]��.�={�eW���oY������1�b���%~�@�*�?0&��1}C��'?��3>�i��?�J�6
,>v�����u�ǎ�N(����ئ�@���ͦ�~=I9��������0�/�����s�����Cl��L���PTA|�u0�ZEbu-�7%a4ڙ|�!�F�W,�0ů0�~��#�f��a��'�p��Sn���w.\x����ͯ��l֚l�)��?���%�.�a[0�:�rW�S'{M>��5y��?9s��#�Ng�V�Z��o~�۷^x�E�IE��
s��խ��shp�֪�1�6Y1��x'��~�����A����.��9p�8�1��JW�Y��c�r4��&�X�=�9F���Oj��s����s���=�<󌫘����ȡ�������<�OB���9��0��D���G�͜9s���5�;����n9s������)V3��M��F�_$DӼc3r]�b�i����}���p]�*����n{<��7�Xr�Fͮ�̥E#^7�n��[9ZKʌ%
�y�<O��bq�����M�z�u��l�o���F�VϘ��dN��m��ZB9E�1Ls�V�PEl�g��9�m��.L,@�nR�'��ko�w�̖��d�$Y��N��Y�2�2��);_�1Fw�01���Z�㴮�ũ���e˖e�I��~�'�R6��Ea�:�C��δS�7��sX�R)�OW�ߣ��[������3�<=�Ѓ�����a��0�D$�E�b�?�R�Bm��F��ߴ�%
UK��8����������k��RƧ>��k_��SN���SNy��]���o������D�*���Ȓ��0&��3�o��V��R��^uC����oe���対��Q�}�����NZ�ti��;�8nqk`j"�)s.I<�5�MǞm+[=6��e�qI�]�,tH�Q������E�_�S�Rؘ*oZ��0Y�S�_�٥���?w���y�G�������s�����b��re�` Ҕ�S��M�M�16��L.� �@nj&���d��"a跿}d��~��Z;�BVG#����Bt�i��p�����?�~�d|���G��bT�������1g�Li�500 �o�m���Z��e�]�p�%�Ă}cS��x�)���'�J��A��f�1T�WZk"������\�믿
�DU���@.{���HED5�u�*�EIh�������ъ�C�}��-�@�R���䮩�b�������A��
�a{{A��_
,&�䁠�	~?����z�>2�E�d�7e��IŜ���*��ۻV�%%�@���(��fh`܊봮p
�$/��v�$�K�'���Hg$ҟ1�j�ƍ���˚��(�0�p���5�؍��0WenL$�\���	�8��c4�1�S��jPK��~;Q�uO8�1�J���h����8���8~����`&�k�U�u�!�>�ĸ)R��c�j���)x=���uK��Vr���I1`";���̶'Al�oܦ���ٔ�k�o$z�By�ιNKJ�LF�h�WM���uG�Ҟg�>��0l�YՊ+�-���O"<�~=��U�o��#�h�Z^�>�c��Sa���cL�X�dQļ�-9�X�x���-�Veܵ� l�^����L���X��Y��Wl�h���s�d�+Y�¤s�� �N;�v2I�Os��78����
è%�d2�f����i{{�@+�;a¸������ř�>��<�(�j2Yq�o)te�\Τ�����~��ex`�6a\|��Z�j���^{�<<[���':����UW]u��>���o_�`��M��	�#�Xj;Ԩ=��pR�@d󛬣ӦN�J���B8�?����p��_�c�׹�;N`>�T$?��{<��*�-�܃|{��C���#���?���i��0C	���8�t&�/7��,�>Dzz�!�7�8�+��leSn�H�:a��$��$:���P(��Ƅ	�Z��(�b�{'�K��
�o�N o8�Ht��cpp�mS��Nr:'�� �JUBMz^�D��&`C�rH�q�R�\.	xk�4@�X��k�x���r�f�Y�(�[�2I��V��'LȎ0:�<��@:)�R�,S�M@�^_�]�1i��Ġ�F��[�ӗFI&%�L�HI��tOE��e���D�1h��1�@�J������iH�#Al ]g$����0��O�t�ϲ�U�'��1,��@L�EO�\�%����	�sM����w7����,@ {ǟ�ST�BJ���}J��3?�,N�s������HH����wS9�����\�s�ąw�YoX���&�a����&?K����D���g����#���)ND?�*�)Su��b�'�3��L�;�ǡW�S����:H���xA�`�a}B��'L�m�N�u�������2i2� ��g��d6�c��	�f�!ʘ)�{ȟ�MaP�Uf��R�n���ɷl�XS�w.��_�f�đ"�Q8F�"z,e��'�I�Q(VM����G����uV��V�R|6Bз
���xD)��a��cC��M��Z���.�X�0�`���Pd?�C��a�:���EB�O�0�8�>����l~J*��j�Sh��3x�[)?��v�ƺ��N	�gx�"^�J�L�c�x`��0�+�O\��:,�׷�I�*Lm��̘�*��e&�����:>�`̵����Z1��e��aa`x�n��i�j���<0$��P��q�S�x�@��d���ab�ۓW�2��	�e�vT�Lc�p�g�͟*g̺�W�L�$�0a\�݋�����|�s)'���Z���d���~z������_�P�^ه�"k!4�����e�[��^`���:`�[5��&ˈ�}�&Fd�S����a��hC�D�k9�m��n�F�U��2�D��,�4��BoQ�^����C_���ڔ�|���O��''c�3V�Cx�s�]{-}����ț+�`����\8���+�h=����++���������|����Ь^�����+_U�}&5^��yU�_8�4�1a�8���y|�������rՊ���N�M}���'?��<�����[�CF�Ȼ�������p/M��5cƋ/�Y]�-E:��(���ul���,5$7cF[��[4���#�X�ݫ�Z�:��k>1����V�~Xd!Ϝ!8��&Q`T*7�s*�T'����a8�N[:AնxU�-vg�R���g	1�ޠ9'��y�rW�^K�Лc��k���J�8�2���yQ*��avEp[~���o��Lyh��2�N+��]��SO>��1���ʹ"/m�N:��N��u���o���z#������&<�|⫞�5��a6���i���cPkPF�[�0l;��e�2�Y���E����~߈�]���Ӱ��(2*�遨�S,v��I��������l�a�2���A4�e�6&[6�Ҵgm�1�0n��?�;�����:u�df���%N��<6��5����AZe�������wڐ�E5��c*�����Yfª8*6�{�:n"#e�3FD���15�f��K���Ղm
�TM}������B���H%Ū�;N��xm�>V�q<�Ib��f�v=2~z��~��j�H{��^s��7�ڊ�������]uH͇�{vY��ӴE^Y<Ł�=�Rۜ ��+�� �5n�7z�7F��l�1�]z�7?������O#�/N��q[��'��s3��&��1���t�)�GFF�����(ӂɏQǣ�l����:r���L;��^s��6yٖ�ڎ���sh��������>Y��Q��m�o��T(l�m�{��]�2�,�a�ෞ�e���J`K�cID7
׍!P뇬��\ެ�N����j��/��y�5p4��>�v=��΁0GE�c�v�1-�@����۳���(�e��ݨ�{�r�Ƌ<�۴׉;0��]��H!��M{6	,����
�A�ӑ����y�в!�R�y
����:'�`k�0e�qVN�6��z8���1���9�C�
a](d�Q�Lo�V*9��08p$3Q��4����<~�i��R���*Q���M�ԫ�O�;�����l+�E��0����5>-q�����.��h�.;�`��`e�ژ[�\�VU�{��S��R�����G$�v�ܝ2�IAy��R/Q���Y�y����e�yU�8�E�De��jmE�&F.\��ڱ���pb'O|�뼉v��7�9���Z��z��[��$�a	�p���K+�Ӯs����p�������P�_O��/�ܗ�A�]Z��E��TIt6�l��l��LhU������������p㭉������yÝ�M%6��TF����ub�H��z�H5w6Kܜx8�z������,����A}�=�LEU*�j��6�9M�"�?���akǕ.�&��}l(�APhR/�G�bA��iȿR�'�=��I�=���UQ�$�A⼍A�!��x�^�F�+ejgkg��D�gH&?�K�O��(*Ih��>?�_���PY�V��o�� N]lɬ��aȵ���R��<d��L�� ������FיS֘`�8>��e
m����2��^�~�}y�u�oh�,�01��L�Q*����ג��S?�bŘC��f�cJ�0���Iq�d�m�R�F��ވ�e���(�����"�%?m���]B�(G :�	�4��g�-O�R?�%B�� �hC�7��,�l҈=F���ұ@�G�
�#0a�g�̚󹙔�����	i�0�6"��X��ux��������ƈ�2F��U=1�R��O]v̧Y�P�;�?�A�d]b5مN&��{;��NN6Es+K�PVd�V��m�_��=�}�T	ҁ\+`�� b6�z����� .'��  T?+=�g�������r)
�a&eD�j��`q�C��D���qX��+�Y`�e�XD8F�O�"-��wl�~Z�6D�2�E��&/�̈́P���N�ya��!6f:�(��Ї�7̒�`H(*�f�XBw- �d�� L�ejc%���b��/%<^�E�����KT��M7vRi96�P����ׂ�����%�ʴ��R�t
�R�qP.�F�؇�7�y&e�GT4�� JF �G�����`����+��,X4~�]���l�͗0M��K�h�&�v��)�����x��L*��>X4C�
;)�^#r�<_���o?��h`�� AVȊZ�#VH����5h"����w"�G�χK�]�Akʒ�p�y,F|�T,f�>��1���+zP�D�C�d��"�L� ���L���X;,ZB_�"�!�m���3��I��2�tA��D�
0�V�b��9EԄA25GQ8sɄ�BJG�� ��e�?�)�J�]�����X"�J��|QF-��.�j���0D$�S>/�
>�7d!Գ(U�l,�0�J�r@��<bšDgRt3�����q�r�M�F�T����[�S��V��;�&%n���6���Ĉ���G��^4yc�Ԉ��6�$���(�6-�\H'�p��P�
�MWēMUb ����WFT$��m=m6>D_/䟞(%���D�Hq9C�|%>#э�rMj��P�91�y���#���{C�Ew
c��"�_���ޘ��|���3R8E�(�.�Cs:\_�|Yej��cXcG
3�5�Dk��^djq����;�R%��0�ݑ(�"!��9��P���'�D�C��W�/�J_��{$�(9���,�G$,�l&�	W?T�b�sX��
y�9e�B�
�iQB��}�ܲ��`��1��Q}O��8�|���(�0�c�F��(W��:5�Zdَbq��WT�v�T}�g��}@/*`G�՛Ĳ4ʊ��Uiu�;p��5C�e��D�	X�����	&��(9��f��p�^�H+�X�HqAc��J��4��v��H�[�8�1��>�d�����G�m�,�S�u'�>b�����BP�q}�R�5SDф�|V���x�.j�#6�M-�#q�Í��F��5�U�]�+�M�/L&(1g�������������X�bs.L)	����(�b7�[�2��B�ն�;��w�S$�Ѱ��~�h�T�,��<�Ta�_�
�{SX����8 n~����7#�,d(�4�h�4ŬS;
[�����xN3���"�E��j�ǉ�9�a��8Ƹn�(pvf��7�T�b���Q�Y�ld)U�PրUi�Y���bd�1��8���x��q�k(=A�%W�.N�9@鸇��6��6�H�~"1_�=\���&�и6a@y��3�\l��&��GyT%42��`�q0ڢ!�`]�b�ITi��xp�0O%�n��[X��Ӵ�G8m�1��q��NciKqb����	c\#VR���@�66��g�����O�� ea�D�(d��q�dL�K�&����/>���b�6s��J�T��UWe #��w�*�v�4d�4e%4N�F��L	���XU뺎��*:1�� g���i�h�9Hy��sfQ��$`�cS��aJ<@�a�邖���%bK�h�ڃ5��5��X�-�s�����#�g�Y�0aq7�{&0 I6N�8�bļ�,Y �f�E�B৞�z�Q��t�OJ�Mg�Ao`����Y��<�ê� ���������Ar��^��!�� ��'mJ����2q���sT�2�@��K����(�-��9�	,,�D��4k�:�<�2�4��I��< �: 8sr���T3�;�c����fnQ���i�[}�e����"B�j���w�b��mJ,V=;�&{�Z�Mִ�@F8�R=�aċ��J�.S�]y~�6f�i������W'7��)S�O��DQ���m�PDQ���xd;���xK��d��A?�d�����+N$J_�(Fù���P��fã;�!q!'��������H�O�Kވ��"T=�JL����
|_&p+�'+,�����aQY��?��3���+�e��,X���O4�ﻶ8�&:�h�$��W�'ɤ���9�M�ޫ�rh�e�c�H��H$�XIq�b#��0qYQo LS+ ߫0����+�H�Xs'^�����e�\Wi9��i���I�E���$M��	8�T�8���F��� �jHWg��Qۜ�C���"��:�ق�Ļ�(mz���ɅŐ%J9��L��e+/0�ϊ<b����	�X(s�1R�g���$FICX1���@�c��,�W���=}T(��*�F�
��,o��� �j�)�0��1�ɫiժ�|BJb� �������R���7�o��Z{� �IT���$�u!6I���Sy�^[��A4��K��1qx�:�9C/K��	ϟbQ�fh�LY�2_�.��:�N���(�#�f�N3����>�Hq�!Kt�(gieSG*C�ę���@,�b�����,�"�&�cK��F����UQe��㇅�Jj-���;�#�Y����W(�1A�9*ȸ)����;h(J�uR��X_�q����wS;�D�h$!oڀs*`�XW�5����l����O��sur&���Rm4�{��,�||��2hwQ��x>X�j��!�'�A��J�T*�y&�
�_�bT�c6�� J��1�'Fb�Xm�#*� /@�����4C^,�x9,V:�[%yRBA��X����	��Z�,k�a�5r�a����]1a���ڌ�tl'A<���iPܘ��}��t"Oղi0.(���q���!$y�E&�
s7q剗��P�]��\�N�_�����N��>d��C�X�*���� �o��&�Ԭ=���YN�<v�I"ǋ�:ZL.�j7j��m1�P��7S�6�S���r9��g&d���Krt�z�-`B>M��i����/1q�
��f��9֮s�Q�aa��FcP�L�����s<ǩ"&�&]�V�C�R3i��Aui�w��$��_�TYl�G�%L��c�e�N�)����}�,> �)��0��z!RO��56QbF�V@��i�1'OE֜ײ������s���ryuX��]_��ꄋ���^���*�;�l۲��>E=QAN[��XD �v����(�ǒ9��9��N	H�CQJ��<���F���	Ew	"�1aDl��R���Y�xc#�Zz�.�]L�Y����{2W�dR��fѐ�c������k�#�ֳh�W��Úc��G��D�&쨋��h=ǈt��j��)��Yc��'ކYa��~����L�U���@S��.3G���8iz%��o�	Wx+QM�O�9��Ma�s! }"�P���	#�,[��\
�T��"�Ֆ���32$Fo����x7S:��f"B#��b���u��>�F�:EA�0 ��u� )����(����U�_N�oX�QJ+��j=d��#��ۈ*�ߘ��U51��ŏ���2J�K�������ʬj��M�I�\�I���F .���zVEW��H]�H�F1��]��j�Ni��u�GM!�
b�/	T�U棸J,
ewF�x/Ԡg�pr�MQ�~���§��8u�W>�H=h(1I�B2��b�a�U�C!���0�8��L��= L=��5��&J�5��G	�N���t�ر������2���c
�K��]�K%)����^���rRH.S�bI��aE�"��Dj�L|�����Ig�ћ$M"V�6��� 55Ľ�Xob<B���3�1�B�u��g�5R�	_j��G#3���&!*xK��c�J4�h����$�@�{_��u���RJD�<�OLlDԌAR�K�B��j#"Smr�)4~.�HGx�i�@L�d�k�i����e����hXE�Òg�@#��"3�֐�`���¶N۰5��z�T>73�HF�s$�������J94����������a�a�cWU�� CgV�-�G�hK����6�c��9'��ǖ�M𼂫h�7�Ok�(C�.�M�Ex�r�)`��TF�4D!A���Ñ2UVL���%�BHEmC�)�J$vMPǰ���ݫج��vA`�á"- Ԃ�fɡV��u�-Pe>�B�x�n.�xf��@e�+(P�;��fJ`"B*��RJ���R�l�&z���@����:J�]�~}E4��E�w��|&U�-��s�Ɏ96D۬�$6��]�la�n��%2U��V��g�d��H��,Ca.BC��f�'p���@R��Vk5�]^ac�K�/�7��4C��" �%b�R1QD.��&���r=��|�8#�l��gR>[sE�Fl���:�9��G�ceu�C�� b-zH�*F���'��6	�3��6��uٮ���H>����QO����OB�tq�H@>��T|�]b�=��Q�[��K	�R���~C�Vt�0)3I�Y���ua+.c4�9��G��H/�Dt$�*��<�5	?�!bn���5��'�X�0�cC�������_]��U]JB��Pu*��'�~�ծ�C���C%*2���i�s�CQ�Ė��W of
KV-Q\-����g��p��@��P5�ee��بD#h`*c��K��Td�P"I<��b��\���馩ce(���U��YA��6�Y�9Y������r�� ��^�\�@�rI�c]Х�����t���|��m�i�	�75�GV<"�m��)R#3�K�xQw�;�-��������L�Hsg̢:9�3R�R�����ry�"��T;��p'^NW)���i�c�!{���w��uk������U��Ux�r�i�P7��c�)��ԙs9)�x��ixs��>�r�5��|�,���bţ0�Pn.[ ��VA
e�Y�dޥ��\�t�]\�N&+DЖM���NTJdY���Di�ζv���g�à��6�_ˇ���*���`�*�%�I�����ja�	cc�.I�x�b�Lg|?z�e�'�7P
������Y9{�fP��3�|ǟ��/�P��)���R�r�H��}팝��K3�6+ǚŮ���]������3�U�pTS�\*נx����R.��b�`�S:;��,xa8|��^@պ'Չ�s�Z�*��(�L�" �2b�gsm�;��5R���4���V���LA���v*R.D晋Ʈ4P*Q���JuO�7��2�<g�#�B*b��զ&��h=�����% `�o�#́�/jh.��57<G�y�L~o��3��3OڃY:@�W=A5�sYތH�Oc�&��A����e�Sɢ�5͞Ӭ��i��i4��#�u��D��5��L�u��a�`������6�������I�:�;�8T��y��������=��C]S
⓱b��������S-ɯ�T��ďA�j�ژ�Qq-�S̩�}�N>VS��w����+��)�E�P�Z�klvQҌ��U���T(�,>P�J�b�O@%v�hM�F��<
m�=����]��󎦽:��������Oh�L�����f*�]s�3��&N���g�C���V3[�@�4�4E�_�5����7���1�{��Ī�ۦS�u�����wҒ����;�F�z����^�ǖ,�߬�:+�(�]G@�Jo{�|�6�[�R���2�˫=��s���A����6��޵�n4�};Z��rzt�2ZSdn6c��F:�s�Ϗ>H��:�FE#Cw?��E^A��b�*9�/eM���;�=�@��	c>�2��$�2LV���cy�tC˱� wb�O5!Y�ev�V��%ϧ.6W�t,q���{�dyfO�z����TH���נR��U����B�$z�L��^��v���o{����_,"�0��2��3��ϡ}�a�Δ��Υ��w.�{�誟�KSXtt�N�s�NL5W�m>辍n[���0K�t�>�h�;�q��4�Ŝ飴]t�r���%T��m;��>w�,�ޟK'��?���h{�]�ɺ��}�mM�DԢ��K��C�jLS�X�o��u1�sR��xuCխ�ݩ��P����Þ����O=K�f�@eF
��TDَ<�q�+��_�N�6�˶���n�1+��n�~��(CCk_�?s<��D��@O/]EUՍ?L;���^T��*Ma֎�co�=EG��m������S[@�ٓ���K�����N#�+g|���O'��jƌ<�Ȁf���`G�&�Ǘ�x��.Ru���}���鵥���DN�j��D�ͫ�D�|��5�)�1���'&�%��8Nb��T�e6��gd�c�Cec'�J��.E�L�WV��j��rJU�>�߼�������މ���V��T���Ot�^�U+ג��A��p31�����=����)8��t��t����>���|���_)�wSG[��Ţg]A/��Y*t�(Up������Bއ����Rɤ���G��ȓ�ߖ�~�`���=w������~�`0my�ӦvRƝFC3�r]�T+�N:R�q��p;���g�a���.��t��С{̡�|��W6�7����>�gr;w��U@�6[=�H$Ш�P�D_Z^e���h����H<��M���T���c&c�-rT_��,>}#���K'���t���oK����CV�2)��E�jm�X"��&�,��;�?��~������_!�}Gr]��̻aV�	�urbjZ�n��g��wn5h�C���}|;�cv�~��g�}j�fg���:���O� /��"Ųf��X`���=g������&������W���<��{������˾y
=�2s�_<NO=��ܮn��Y9�E��{eo?��S%9{���K˗	G�u�)R��ηK��g_x���v&��L�
�$�}�e�R�*	��;Q�vC�j�nc�4GUhA����C<�JG�y�$�ꬿ1�Jƍ���Nk�B��O��=_��6Ņ�*��zY�ɰY����>�	H������}����NL�_�yz�Q�Ko���A��LA�TI�R��葕颊��H�m����u}�����L�;�$č�zm�z�dQ�Γ_���ZCKW������f�B\b��������VV�}�ܛh���л�K��>��g���C=���)}}��Nz�C�C},��R��M�*���YJg34X,��`�:��"+�[gp�	�(�E�P�W�!�C�FO��=�Di�����,�H�(���[_i�[@���]�3R���VO�
�%��03���̲1i�tɝ:�V+���W�>���nt����1�?�[j�兒�5Xe��k�f��YNէ뮿��z�I4�Z��2)F��*��7�G~��t�G����ffS-T�.L�[W&�Jp���8)�'�*�*�f3a9y���ӭ�Wҭ����oٖ.:k�y��韮�9��uLgQӖ�� �M݆*}EVZۉi� @�V�؄-I�:9<�+�XgE<�fn���W��Т[��ſj8B$k�u�*cH삂��m)���@"k,e������g!,��_<a*�'��)��&"nqKN��e%U1���z�CA�ewz:���􁃷�SNؙ~��+R�=9�٬@�C��U�y����֮RT��>�@��˯��5��5D{�-��c��S{�@��O�7{6E�L9�(Y)��&��,[E�j/�Cm�5[(��@Zߚ54���?��O=F=����N�V3Kx�W��mK��so�颧�(W���#=PD�ݿ{�RLxq�� /W���1��L$�C>����pB1�"��L����R�0��4
.j�b��0b�{A���oF�['�W"8�並�*�@$�t2L �����L�G�Iz�C��R���H����|�?[����˶��7<E�|��t�GХW�GS�fP=����Ot�ns�c����DԻf�,����=w1��'�0�X�L�MW��t������s��ޗ�^�mfmO;��AW^�$�i�R>}3�d�Q-����T��9�O���Y;����h�w��I䱂�ڒ?S�����hG�W��˄m�ѿ�F��mK��z˜����>Ms�sz�M�����WXL�ie����X� bf��0'AV�ҋ�fPcˌ���d$Y=*4���*a�t<%��a��.�k)�16s5�6ݏ�S����$)EGU��zN�i� ѫ��t2�~z
=����f��LTO�iy碷�n��l.�؆�eJ�w�@�����
�|�4�f�c[*��'���_��=�2��N�ryz�%t��K���^:�sD4�ġ��Ѳ���A��
���Y})��ζ.�f���f���c��N9r�cޮ��S�_K�_��D����,�"Χ�^r}����C����'�f�r��k��w>Jv���c�;OO� Zœ�����S�4"�ď�RcV����ƪ4�I&���^(d�ш�*���!�	����F�%E	�3�S����.��`
T�M��s�J6���`��ѓ���w/b{{;�U�6���x�T������28eZ7[Lrn���֣~���L������`����g��B��V�C�C����=�)���W�be�����P��K��U�εI���`���^���>��{�k�j�nz`�tσ��D��NQ�Q��]X5�K��k��ϟ��n7���*��<�X2 �e����^��K^�+���ɢ�g_�;R ��JRyQx�(��.����+�N2O�hbH��e������p�&����g�~A�L���� �����S�PQWVP���uH�j�/	�>@	Hf��w���Q�!h�Fqp�P��FTc�5t;�$!��i�WA
CPS����)TD�8+���`_ޜ���b�L��,6��J	'B�ӻ����_���i;�[G���HY�q2�C�mn�#P��$�XJO�#��k,G>����p�Ä���!��ܬ�d �{K��b�l��3V����4x(�b�O���aB��Gg�t����@��q�p��o�v/�k"�
�S���ME9�5/}_`.���B��À	�C�'9]"�,S����P�[ .*�,-m
���*�WbK()m���A�=�m�+b�s��B`{��Ҩ�㤔R͛�+�F�g?	3�����������
Ѻ��<�X�%��B(=���ʉba�l�j�l]��a����*.p�=c���Y�'&VR�-䚘�n�
,���_�V�RA�H}2�GUAccI Nc!��U��G�e��J@��7�AJ?M�O�@���T=T�A��T
EN|i!)�Qc��P7(.����Cĕ)�{2�Ȗ������n��Mq/��#�%a��s1���"���b��(�^�RU��������� ��!PB�-��,Sk�MJ��!�rb�5' ��p�T�J����Zj����G�A[���yҗ�?���QT�ut5�WY|�'�<��/�k;��0�y1@��U�S���wL��NDo9a[�п��yA�@��*a9�eE�/R��Q����X�6�t"g�)Ś���V��/�`��'R�l$ʲI�Y^ &D�!@8 Ѡ{uʲ�$ռX
Jy���l��5\�y���8�R@N��8�9(Ub��3�V����0��t�s�
��d�mR����8�XԘn�P��V��51E�Y�x�� ��͵���<�����T
]Ή��pe]��]pٔ�P�֕ �X<�K���<���(
�b���yUI�����C� 5��U���	`�+tba��	��v�R�+��,��eQ���	��h��I��@�����ErA�<�j��rA<ӑT��-&$p+�l�.��M: �D.��1� ���LmF�C���!��݉�`���	��@8�ͬޯ�s�r��t@2T��@O��a�5 �
O�*�T����e3қb�R~X1��@2oul��\>��t#I�,y�A��٬bV�PJ���׵�(��6{FG�8Y9ˣ�W�P��*�_���f҂R
�jC�h� ����8�N�ιT���IʋfI�;X�S`�Pz�E�{��L&(xUQ|%��*W� !@�\p� �w6!�)����s1,0�[&B�yl+�,����Tx��[$Y�!0���y}͛
L)����!g�n������,:@U�O�*}+�//�bsHǄ��e̛��k�G���*��<Wg:M�>�� R����gB˸!�X'q��4��%�mTS�@w|B�^�s]�H}Op|��v�ڶ��(�Tc=��=��1J��1���U#��+7^I�Dk���$`(]@C��A$�
�w4��mw��Ա��T\�Q�*$������釩��Ս�0�+T�.��U�V�-�l!̢]�؎��4Q! .^�s��O�-�5��x?��TH�*u�G���z�#s�&;�N����̳V�����]�C/>��'���ST�~K圲|ϰ�8F5u}��#p�}h��?C%t(w��D�c"��x���??I�������v�K���!uN��5P��/���?w!��n�i�������A�o���@���g~��e�����(�0XT��-�4��L&G�����IauP���l�y�!�A�'�v�9��y���
��{���B��N�QřT�'�レW������_,�c����\CJ&�L�Pl��#^�iوf�;�v�1�Y�R��k��9�)���Eǭ��AO,롔W!�S��<s�|�u���\L��wo:e���5m�A�ʞ�,��3Xl�T�n��b���s��l���e��0���Ru�������fNTa�H�/b��h�DA.27~�5t�od�X�����'}�bS�3"~�'��1�5�E��\���6D�n,09'@[&պ
� �D4��giv;��� �Ѽ�	�w�芹�O!��Q[.m�������󑥓yP#�9�\�)Lp]i���*���7|D)E�;�i�	������+�E��iR��Y�E
���H~2���x���# i*�ZET{����M{��Ւ������b���b��כ��� n���q!��q�c�YA.�/�k���^#�Q#ҡt�cBj��F���*K��|�����pC�Ft���kؔ�H꧅��}��iC�e�uO��@�fٌ�E�2��{6��rq���4���3a��|���AJB�p �ԅ�&f�_3���&I���9�p�C�ur"#V�Z�� rB���$B�H�M�	���TX������%׍'u�F=P�bCu0lG5�&�R�R�M�+����q��|�8Pu� f��bԓ����F!:D��y�9N�)����
U44�k���5���yD��bh��-�_��÷�z��Q���~ �lE�ե�)C&�H7��m 6���cH G��(�v��L���-~~P$��R�����n�@��sǺ�f$VNzv�=���4t���2Y�W ��#
!kZ�����bV��L�)1W�r�4BK����gJ��##����瘽{��=� _��-���T�3y$���`H?�x�j]�d�\Z���J<��T�*�L�_I���t.��1p�2��=ߴ.�y����etKJ���{�:�M�Yʁ��߈Ԏ	<ޤf&�� l�*���}�ڵ�7����F��]�d@6By��,�8#�k8�$0��,�\I�'�(p�pU�$����K�Z�|���Hm8E)J�d�Rg�@�#I@B<:���T�"!vd���ä��@�Ռ���
C����J ��b*M�:��T�@E��GWrz-d��򘉠�x�̭`���)I 5?���Q�IٮqA��[8�Ⰱw�y'-^t�,8F6�j�~��E����˧�$�9m]$o��p�.^�.���
���:f ��iB�C�It���ZU�P`�H�_��T𹧞x�.|�/��N�J��}dQxA+v�WgQ�1�\ fE� .��"�^��sK�H�ܼ��H&rTsa$U�	�b
��z��]Ya1���Ɛ1\�UED#���(�?��ZJ�C��tEUX>lt�d��M��\P³&Y�9o�����5��%�!<�._Nk�RcS���q�r͆	
�){���]��c7Q�g��Q����^~��[Ջ��\%��~�4.��F,7|��R!2��¢�� �4ܲe�؊,�e��9� �NA�����i�+�C�T�PA�j|(�lGC�����ء����]R0=f��w��(��দ����a��Ǥ�[�,��T�$�Wzı���֧�s(�h�ƕ{`�c�ch}e�S���/7���C÷�:�&i!jd#`%�I}��l"�憱�!l|����7��-uC��b�I)�O)g���M��i�?��u95�>r�x��-�v7gش���t�q�aȦ&!p)0N� 7 ��=G7߷f8�~�ah�/8�'�8���~U��P}\��bC��J`Ѫ�}t��h]
i��n�f6,�&|�F�HQ2�lwY�jU60�\uBI���.RM[�H��}�D̤R���e��ͷO^�̵f�1��IZ����{:�3Ho�с>(���@�MD�noXA��'=�M�8<GC+¢�e�&�,4�Q��U,�()����d�|H��@�tD�F&Y�h���EJƽ./)nR)P��zS:Gi���T���b���+�F�
$��G%"{�j5N�p�X�G�ԼF^/f�����hː,r�g$'�AZ�l���=4T_5�u'�l���9�b%�ћ,�cP��O��zC)��q��M�Xx-�H��b��*�I\+�8,5��~*��V�VR�]B�Y�YI4�~����'8ҏ�DY�.����DJ���N=���L��Xz$l]m*563�UJ���aqE��d��6�q�Z��78�*����5�&�����Ł�:�(D��'�o�������:����A(�X��$��֩���br;�5G��i�u�HS�DFb�V�+)�I!�ULE\|r�tbQ�j�XR�Η�R��A���]R����|n�\�kl�jQ� wx�MK��_���F�"��Hİ�qZ�L]K'V�U~���|�:���0��Oƨ�����olA��S�E�tm��X�%f2D�IM�XNw�X���0�D�$AB�����7)
&iAb͑٤�5�X�r�H�q�J�׎�EL#=.ɻj��O<��-BE�5�'�
bڊ�%��F����b��0�M��#H8���/z2�eS�8N乮5ּß3�T��M;���Z8ĉ&@�@b�(����Nn�7^b=ڿ�|�GҬ���$��\�x	Qp������Es&���Yqn�|�5"�r�?#J��@�,�z[��@�Z
*a(΀^1D|F{mEq�_ƺy!� Z�|����4�Q��x��{��ـ��3}M�\�ډ���xƖԝ�8@�eDB�]�E��<)&�>�&�$Wץt:K�(%#���$nr��f?�'M����:�ǆ�a�s���~�+�r��ZO&�����M����D4��������f�~mD�%lisyx>�k8I�ў�X1��F��9#)�/(�f#"�ՒI��A��-5��X��5���ؔ��:I��Γ�=*b8!۳��L����bSߔX�/��0󖕇|�~뇆����8(3W~*�qC�S������3����[h��o�nh�=)��?D_}�K�S��Bۡ2���+V�A�5���[��W.ن����UOc �3���W �4��j������ت�$��_mW���'($g�hY��y�9��o"t����R,�u5m���l��wI��ύ�(��I�l)t�����I�H��:�ee�����q��rP$y5���>��8C!�%�,�7ְ�8P��Ke�cO���/^F�G�Uy���"�,�f�T���}������]��Im!I�������G�%UC�Ԙ �� �y1~��o�k��{2kub&�����Z�i��ZV��q.}���yC��	tP�L��� ذ�.ʼ���~�a����ӨR.�:&�~U�8W��+#e��������c`�D�2�Q�X���^we���G��:���t>h6^"�����3im� �ӷ/��D~����R;Rj�1a�wHFv��M��CC�(P��q��d��j&�Y*JP-A��A2U�����Te"�{��l�[ �:R�q�LS��-rR����s(䲴��QP#_��
^�z/�S
4��ç^�fT�&C�
b�/�@��K锋lR�yS�  �Ђ
���󔚳-}���h�\�t�cD�+�ӓ0�}O�@��8ڼq�.�o(�d�am����>�)ʙ��³	�#P�}�Ȧ]�Y�:����ԙ�P S@�i��zdk����#���qX%�+�@R����X��)}D�TֽPp��ՙ}cC0$�� �a�^�veG*�!kCu���Q�>M���-1� bº�<٬
�#��Uw�$�\E 4\�m�.p����!�P�sF2S�l��<�"��Yǔ؋�Ĉ���r֘;����$5Da�tB%j��d��=�|���I-H��*�-�n�z[D�� �Y���C�ֆE&�Z�����5�Ni��@�!pB�ZC74�z'	ϛ�*��V�T\��>�S
3�UA���
��)���Y� �am:���E6�Do�q�8l ,�i�]��a��, �ZI-	K�X��Ѵ]�y��{�U?�5�c�*/�a��Î��c	9�ir�4���(#�<�J�R���YY&B�9+�U�k�G��7�j(�r�(џ�������6�"T��+��"E��G�H����%�2HE$�7�xk���6`"o�0�[#ͺ9���2y)��0t��ʴ�Z�x����](�	������e)�e�Hl�Ʈ '��,VA
��Ϙɦ��pr �N��&�j| IP|� �C����AҸ�HR�IԵ�@��㴊^�VH��H� 3pS�/�X��r��{rr$����h�R~/a��H����\L[~5T:�'�A�JAL�ؒ�&X]Et�W���`��A;ɿ1�x� �Κi`�jŊ���{�[�U��
;�*Wu��PMGRC+ �(�p�>�
"���lT�\L�- ���%�D��n�s���\'���s��ϩSU�T5��}��+v�s�^{�9�s��? 6P���{������j4e
�� Gd��zm��tݼn�t���[@�.i)q6�0R��ܥ���	�Mم#m"�@�:+^C�xl����2!�����ma̜����J�,`,GS"��5� �\l����u��! W�\B�0�e�}"�p$���1HR�E�a�vN������H��S�o�R�A�K���d��bcЛ!��������إ�d����5,e=٫m��z\�ְ^_%��5�l-\���We�#|����O��2añz�\�
�S��p���VD��J�b;���v�u1�F5�,���J>�wi�BS�f�X��!���u�^(�U��He!�q�\�\����b�¡�߹J�m�AD����H�n4����v�Fq]��~o���6F��P�����������gMT~��螰{=�v>H{i�����{䋍��)<��/�6�d.�OCTkl�0�����g��U��}��U�Zް׌l`e����'�"��ᨅ�v�x�-\�l����#+�	����Ae���ρ�!�(Ҧ�����p���H桫;�R�nӊv��d�<�����L���+���%�XT����%?��=J�=+�<�K���I�F'�k/+�v�U��9��6?��}�Zg�*��[Q`�La�XeA;`O/V���U�;*yttȩ�q�/]!��U�"���tG��/Z ��@&BW�3��|9���Q�B_�F�-��X�Ќid�������2,O�.�!w�K�A�X]bd�Kaf#�ʀR��!�B*цQ6��q��ܴ0 t��U�A�:A�� �fcQX4�����)pH6Q���Y���y�]��i��.Ϣ��f* �nL-�v�%�]��ZMVJ����T�����l�,.LmC�,�'wQI��FS��_�8c��^Vny�Y�RL�GDAe�i5�5�W����p�0ϲ�<)̂���`��et��� 4J�><�1,	�6��)Ѐ��+>0s,���B�Y�m:AQuq��w��yV�oҎ�»i��*�`�vE0��'�ob�@����+-����"��L����H:F�_�"��mjC��\�{[�	��s=j�LG�!�BZx�z��8IՅ����.���Պ�]T��Ŭ9�ՙ��υ�}&����j��)�s��	(��UXw ��yMթ���؁μ�,i��PP���16���Za��U���X��������+���M]����(�o�pK�z_8�Z(åp�8<2��ƁұN4'{�_��)��ܒ��z��͒.�B��#S-I}��al��|�ν�

�͊��/8_�H[��.��>�,qU,��k7�3�Z��k�l�؄2�`H[�B��,k��y��T5AE@_'���I��m����	5zi��Н�Y1��3#
���<��f�F�}�;��L�����8�ź
8��C�ݑ��pz�b'���Zp���3o���[���1*����<F����-\f�}/�@εF%�Mb#� uc��}X��ݷ
�.D`5!�������G�\~�:��8�q���P�h�k5�.t�[>4��Ѣ��otR�s�	P��깎� {1���s_�,1NRY�s�ե�8���u� 3��֪����.SF���zt=�%*"v��PP�{�Ư(��5qWݼs$a�,集
,�P!��K�ّlKo����4��Y�gӧ�Wg���K����T>�3~|R~�ޫ��0�Q��XN ��˂�Gi�-97ͱ[h�U���`ߏ�j�	DY]f0>�&�XPL���\�AI�� ��|�C�|�v�Y .T�{�����[��Z�w���pж������5p��l��✹��Zs�9,r��!g|�
��7v�T�q�[H<�׀%�Giuu��PL(�TG�vY1�tn�,׶ �5w6�-1��q��~���7�n�=A���]�ɰ�%�UQL��?��ی[��������D���wcY��E7e�n�Ge��TaƲ�쮪t����:C6��J5hf�N5��@�����ӻ��j#4�5LF�wzd�w��r�Li�̭���`"�{鉱��(\ř~6T?�` ���**�V?��ĥ:�X%k q:kU�;}ͼ�Z������HS����}ZGr��!Υh�u�l�$YҬ%� �l��F�DE"���
��L.��X���@�x`�af���<�>�h����`�ff?�����A6t�^U�$
,:�e���a&x9L���bh�
��/�Ԡ��c�2���:�Y�`A�9��/��$a��硆l#n�2*�r��瞑ZX Q��QW�Y>�<�`�A�nQ�UH=Gܥ#��Q3bx�:��I���*�D��պL�����D���P�N�-��6�j�g����b\.��ws��2]�x�C�p�D�����C�G��%��pp�v^�8�yO�7��
0�la�]���!��Z��0C�x�WG�P���D�I��>��a%0��Tpa6���j:�қ���<�s/C�3��x���J�|�g�>s�΁!�C��~���}"��� u�-�)f0��`��X�1V3EH^W���Şu���ݕa��IbB��w�^�EB8��P�6ѐ��;�W�D�z��$�A72�@4Ks�z�|my�����Jn���%�����!�4!���WZ8(��iny�^�D�ZD���Yw���u����JS�� !�U"cĬ+mm�.��R	�
J
gZd��-3r
e4�4
�g�<!q���,���0�%.��dlTDd4���P����������P3�)Q�������j��������/w�F��6��?��r���b�G�%��l����`K$�I��eW�����\��7������������!�|;�>�v_���|�&.���!AA̼�l�O���%z$ϥ;L�Zv��t�V	���KQg�,�(��T
�\̾�y���~#�'�Z.[��W}6m�6�sM˻ ]
;+�@��
�}��f�9�f�G�j��1&�A���
4>�:�>�tSm�^q�B7+u��^p�mw�o��>Te�eH_5u�,^���zo�B(�bb���;����mh$�)4-�܋g�}�F�T�$*.��ۡN�W��-���,��.��Y�*v�y�\��
9��ݻ8ğ���0-����i#̓d6d�YS��Q�Q��w�43T��<-�{V�x���"DY�����OGd�q�0`�42���������Q4����ް��~������ŉU�m� ��pWDJ�ߎ٪��\U� 5:&�����T�a&i�Ҙ
/��̶���z�E�����~b4��/�E�Wg�R)_�ٛ+���5�C�7�ό�شc
�c&C�����Ǚ�6�s�U�E���2�-���aT��k(GU����'��T��F�`�o|��ȿ�Ux$3\�9&J劓����>�pn�]�	ga�1D ���9��N,��	>�8��HW��*�}�,�|�`��W�m�O�Xl��3 �bע��}�f�r���+�0�@��͊,L����{r�K2�K ��c���i1";�i����-/C�N�ZB���-9�d]Qrj�2�9N�&�H��̊���=�ϵ�4W��X+�G���0%�ݨO�{�n�v��6��#�in��$��5(
�?r���쇻H���E���1T>���Ԙ,�����6�g]!��}t������|O���Υ,�!��xJ-@5�"�*ɮ�z�+���'�S0ږ�΁½$��՛.f�3���"{C��I�B�}�>�X��ϋ��`h�ܣ��E�
�/h0�р��QXÒ,��K_�2[�>h�7�Uq�D[���l4�:�Z���ܠ�!F(�B����=����7��n��;�F����zzSvZ����fw���M���0L�T���Ȫ�#K���j�3��f��v��ڝ��wYp�G

6��c	� ��7d����^WR��2�hN͡GHC�����E0,��ʼ�US��(������5F�סU��R�)�
�X���*e�(_N�b�0f4.�>���Tm�HIIe���Нi^��M��&[���ɟך��~�\��w�Ei-��i��k���Sb�,n�<���F�sT���w��-�$�f1��s��4 �tM�Rr��b$uW����*��|��iw-���.�Ϋ�
��&��:53'�`�p2u�%#�!������ה��P���ke`�Kj�2��n����a�C��,�%�J
p�!u�W��P�$tY[U �Hw>^�cÓ������0�B�M�o�>	.�1��ݾO��!`� �1L�P�0\ڨ��r��ah�AUl"�ϒj�v�u1ִ��`=G/Z��f�����0�0��K�Q#�Q�ѓ�C��@��}:�=b��	�Y��\f+�Wt:��0�PC4좑�P4�p�Tu����,��@p͚�ϑ���a��r�n�|j�Vj^�>�X]0��T�;	]��ik����;�:�p9�xB�qu��C�'�Da�պ�0FCw�裨�������	��x%6B��ev Z�뿎Żn�x	��>tn��y��X諺U�0��ynGq����ð�I1��;o�[���Z��j�Lե�s,�9}|�C�ð�F��*�{�s�Q�j���7X������׿���[s<[<�w�󝘒3T�?�Y6�Q��� W���݊~�t��#?����)���(\8��' �b�Z���s�v�DMͤ>��3�)�q�h�5�F]��p�5�B[dՄ�zwӒ�#c�ӊqt_KTv�O��v��ۀ� 6��\O����-c<�5aF�GVm
�[�c4b�E_��W��K�ߊ>P�G��=���W�0�5��nY���Pc�I�d�k�{�]s�w5��[���'?����"��������ǩ��0+��6Q�fk���5�a�qQ��%�&8��c!�o��@	N�1I'!/W��(lyc�Q�<K���^'=68H�qA�B~���0���ep�
d�Պ%ȝ!�X>��i	�Iu	��2����G����MEgD�g�A%�L���#�b('�,?�C�x\oԔ[�%o�LfM/��g�NL$�W� o����F�F-W��A����z�P�����:�CW8��'�l��ԁ��p[��ŧ��1��,7�f>W���J��J0a��i�c0_��p�9\3h`1w2��/��X��Ɛ��!�e������G�����͉�E���\�z<��;��� Y�2L����<`3��+��+]ݴ��n�s1~Vj&���BSs�D:���� ��!��"��D{Ք���+y�ۑ�H��X�4PF��A^X'��OF�$�(���9��rNj�ɲF��^���a�,L��>sJ�\%>�6���H�Pj+~�J��-\J8��s�*�d*����!{lt���$T��d,�K�����v&�n��R�Z."�Mt?X����\^&���5bEV��H��G�T/#�ˣ�O��c<��h�m�-��lsЩ,�
|
��N}��qҞ�\V��F-�v������F�%,C)�j+���tz_�s����E��=��R�j�0S�si��l�[4��eyc?���Zv�%y����l�0i�\�Y%����p�ى��^��uW&���3����m4�Se4d��j��r��\�ء����׮���������XHá��W��9��r�3b�u�7~@ꈀ��U�s�p����i��3�z-���\�F%����Hܢ�(�W�ԹID���$0ʊ�0�Ct�*6?c6�V?jq�����䮖�ԁ��y�P{�QrG儮f5O�jy�8?����劣�cC|ٟ�/��V��u��:�YK�4���p�d������B��b�����zf���>��3�׺������h�lҠ^��f�S���*Vh��C]dj���!,,�Ccj��h�kDXL�$�z��=�Z�J[	w�K��P���]��13�p�uX8�X,���+wlP��`�Z���X�xbT�:b���a�bLD �a��'�@ֶ�z��6Xոb|wĀ'�wsfN�K�b����Q�k?�#�[��[��.�$��F�k���Z��`�#�� �O��fU�b�V����O��d��M8���H��X٢���f�J�#N��B�ZeZ���μ�"T�ieVL���Q�0��=�����D��AY%cS��A��P�S�qR��5�ﰿ�ܪ�iH�=�B��3��W��/*�͋�ُ{���oV��[�0�q'6nݩU�D�ٲu;��E�sF�Q��Ë��Cp��3l�n����a�����X�N��R��q�]D�]¶3��h�u5<��޽���_�+x���e�y�h9^f[b��p�w���}����s�05C(��QmlG_��bs�Y��Z35�����>Pv"c�����������`����'5�5k���{�`��p�����?���6�U�%.�d��G�.QwX��*��X,����{�w����;о�غ�Q�u�` ڦ֘B��]|�Y$b�(~W	}ߌS�$�50��*K�h��٬e��Cr�����2�ۮ�]����ڌj��ޔ܁ͧ��FA��p�9���5�Hs��o��G����5��3�}݀Ab-�A�2����$���G�	Z+���$#-3��:VP�1��e����p��ؼ�j�ɹ��[?�]7|��kO�G��AqMOd�dh57b4*�I2J���>����<Įͳ�=�sӗ����T,C;�Y��J��pB��R�2Nr��w��'9*��u;�VU��,�b����[����_��?v1���/��s����7݂g=���W��٭h���Q�"m3�?{��>�q�>�t��s������K.C�9����7��g0���	�ic�Қ�5E��2>��A�&j��_��C{P���/an�"��~��ֿ(d�7?��8��]hGm��]���|�tӍx��~oz�_cq� j�Z�6��uo§>�y�&��A��K�?7\w5��18���\`���5��?�J}Sr|՚-9b3@1Av�`�� �W1"7l���� ��!->|׷p�Eg���y��/�Қִ:�t��E�X.��|����g?oy�[�`�E(^����شq3Z�SZ�ڜe��H=��/�?f�؉�����'cnF��Զ# ����*|��r]'2V�DO�k���o�͠ڌ�_X@�x'���g]�{��y0���w���e�k
��n���]���/�Kq������=�T��]BF�(ǵ�݋G���q�/�<���{ދl����3P��&�����2�t�B�qJc��`�D-�`���H�:6NGX�� �q��.�K���g>K������s�t�mk�c�y��/~��睳K���DTd�%w�w�Kv����ڨ0'��?�����w�̳��\�T�2^8s�8Y{�sU��`����LqcZ���b� ُ��{p��b3�G苇��g�� ���û���Ӵ%!��}"�u�%���M
�Y"m'�V�bW�$B� ��oԞbc�� �s����P�R"m{��;w�x�ەl�k����S���%�r�
�9R]"!�r4���B6w�zأ���R�h�����g?_��y����(GG[<����#��h��Zo�,��7ߌ��/ğ��r�v`������.�o�q0���t�����(���O�g9����z����V{	ƂR8LgZ�J��$b~�0zK��P�g��x��]�L�,݃�-m���5���bt�\������'�u�����u�1.����܅�/����w-�E��"]v)�Ze��{�ޡ6G/_@%l�ݚFczڪ�
�q0��p�j���ˑ��T�kR[(敫�����()z�ƬW�<q��m$�k�����eg�Ш��s�]���06��!�i�u��WkX��Y.���L��&��A4�����P������J�(B�6i[$V�	1E8�t�be��)�q��`�E���#�*c�cܒ�5�$�CZhWW�;�f��ލ����E�,uPW$�PqA���/�u�zl<m¦�(DX���%��7��s7����/x�s18�u"7�e�aϡ�\o�μ�B�$�+y�0D��-��}# >ec��?J\9��g�UD�'Y�Ѱ��[eV�(����]���n?�n�zK["?����^�R4ڄ���h��7�WA�A������mÇ�}�d]<���m��#��;�ȽL#I����\õ�f��1�qq�b�e�Ȫ'đq�S��e#
-'�&J�a˔aHvj��g:[����}�k_����0]5\�/|�x��_����y�FYO���r�x�uZַ{�yj�Fu�N�眿��G�i���_Q��T_��7�8W�����g���v�]=��>�1�3
�Z8���:��� @俉��N~��eiQ^����p|�<��/~/{�+133��7!�E����q;�6o¥��_��c登��Ba'N;k#��m��v��>�ױ��a|�S�ö��������e(d�J+�I��G�����`gxnu#�	5�Ɏ�e���v��ߋ��r4E��[/����ϨF)~��/Ŗٍ����1,�J���n�NO�׾�5ر�\����]���ۍ١�nD�~fozǻ�ܼw��JK�Ȼ�� ��Ѫ�(`�A/�k���S��GqD�y9&k��"�j�H�4���+�'#L�7`�����;���/���z�4ds��֔�]�y�]������w�@��x�k_���J\s�wp���ik�p�G��FP��W�Vi.��_F�ލC��8�ZX�%p��0�v{�5�������\�uō���1فn�������ô���Qco�/�S����'��ϿQ]w�q'.<{7�K�8�� z����`��ͨ�ut�4��׿	O��_��7ށ3�:��y�D��0}�#EK��Ae��ulk�9x�
�D�j�����<�1t�X�I�d\�h��H�6@��j��im
�� ������c�;����o��ضm�x5�Om�:��--���o{3�x�p�m7�='�h��7s@�t�{��:bx��<	�偅:w]k@� 'S�ud�+?��p��eK`t�߭�1Ҹ��a_Q/&C7_AI���`��D��k�����x�{��v��~���Yt�0�f��3ӱ����Y�{!n�I\ӊh��s�c��qסEl:�t����	P�q��%�fS6���qJc��H:�Ө����,����f0�]�<Ksg��o|O;7�3�M�v�=�ᰂf��5���-"B$.�]`j�N��&�/��K�}K=��y�r�M�v���cv�,���xg����5�c��5����\]j����w{#eW&U����&"1,j lv�y�
9fq���;��$^���?y�><�<l&���{R&�O~�����3p��O��܅�hl�s-q���s=�l٩�}ڋ�	z\���Z��4F9ֲ˖�/�-���,�k�Ĩl6�O�Z^�����*GKv���3 ���WP,����@ܞ��{2�a"����1�s0
U+hLoD� ��c|Э�9�S��uO�3������7p������3���r�lFD�򤯋��"dX��޲i��,�gsl>�ǔc���3v*��2 ��X�{ϋ�*
�6�y�<߄F}�V�Ȉ��+\�^�XԒ�+%��/��������ʗ}�(?o�]����0��ϗ=k�3����_�&����6�1d�;2�sH���/���*Xw�~o���=�����(ĳ47���DUm�D���"�۷Ga��6�R6��&H�@N�K���+b����#l��F0�˄�V�T��KCT�R萄�2�U��A�I�	p�zc��5A-٧�Ȗ�$�F�7��n_d�:��~��ZQa�t�K4�������>��(�jJ�C�"����/�ǣ�0bT: �щ�\���ص+��D���*��ـ��H���I�����7��P�C����C�za)[�g]`�r2�d60E2IZj(��J� M�תW:���"�-��"5Ɔ����x��/�Q:�S�a�G5R8�@��=T�M�1%�y6BK��c�F�#�r�Qd]�,C>��>Eg��{�������6�/�}�����/���G��Ncl�4/�**�S����ˏ��WǄ7b�µBy�	@�b��exGUyXe$�L���=Z��]���I�Mrg,.Á�M�،�j����>��.
C�ue��|��#�+]��/�4x��j\��u4�R<;;�o�TQ�Q�D�<*Z󡛉��T�+���Mm�X		Gz�Xo�E�J��.��A4k#�q�5�֌l�)�S��ƍ;Ā��� ��FT�<�ZA���9����)[i$���/D����&5rZ�w���]FH��MA*�̣��Z���r�X��?F-��lT��zA�ץ��/�m��a,�P�_�M�D&m�hRt��V�����J�ԇ�X_�Z�X���b�|bG��x��P�Ȇr��9��W�`�T�f�`�Ar�C�؆UӟS��)*������u
`_�YZɽ��ĕO���y�]����k��M�[�Z�i��}����l�09�Z=2$�9wؖuQY}�Y�c閁���$\��f��5��O�d�G���Z�v�7�'�v
�?&�X��A*$�_�y�AODbńp������O��Kx��_߱(�p�Q���(�INdc�yi�W��rqn�E-o��D�[�LP1Ru�Yjb.�t������h�4yds��q��ɳ��e���Q��_w��tu���������e�P��5]�7��H��}��nwZ6�A;��Lz)���פ1��8��l�-7�X����UQ�Ia |�%#��%��[W�����w�H�g�`<�q�Rڬ�R:M���ڥ0U��3���v�$�i��d	?w�&�ɯ���'��h;�R���1��͡��.��9�q(����兯����(0q�x�=r(�99Y��T��UqS�*C4�yZ�-ٳE����!R[��[ɺ����}���B��[�Tɠ0H;x�/�,^�a��)Ɲb�.����Rɳ��A)�(�(C�Q�VQ8�l^����pUk.�X�?���\��1�s n���&�ŗK���h�t�f�,D�<��Ύ�J�a�:���@��N!J0�D-)�6�f3E�S�c�&�&���Xψ���������í�G��ޗRO��yZ����EV
ő¡~N8QT8\,��OP���8(I�u.�ٝ��3���P��CA�-1[�㮽�`��I�N4�Q(dÑ�%y�G��h]�@,���᠇��ѣG�e��*�M�L�b^�h�t`�C��nCv�?p�_J8]�I��t3���[������(nc0�x�K��)W�=��Z�'�����:�R��>�w\�s�>�3-�� ���t���Ck�9��[ŧ�������.<ː�s{��+�5�������� �p���D ��j,
�+RGD��5r�O$Z�P�d,��TwǎJ�kj?w<���f�zL�<�w־�Ȁ���نc�{����9d��0�o�:���hk;��:��b#M�30X����VÊ�V�Xa���jk��П@���1+36�����%����-�Xh����;�/�e��j<��y*����V������?O��<q��cœ��P�{����=yc��f|��+��>�7��qC�,�s��H�i<��+����~���ص�¯�ʯ�[�:���:���'xȣ��o���n>�#�UG�%qp�R��e
c+K����Dt���Rz1ˇ�'z�/�Y�Jǡ����!F�mPJl�J�`k�����}����'��]g?Y��D���*�E1�?�����{j�i12E�U�8q��5���,��*�w/�Z�`V���3��*�ܳZ2eZ��D
��]���V6�S̠��`wP���	m����n���,�XJ��p�Vh��(����Đ.;���O:9�bY�O��E�#N�"#5�*t�����^���)��F��"�F�C�5�YNG.�T� �P������J�(,�c�M�h�,�6�l~c�3ч�">��(I��,O2��������'��ۂ�X��o������0l�m����>�)�+[��8<�(Z���D�b?Zn~Z
�k�5��Ȯ+���G�o&��z"͙��h�b����C�s�u�Fb\�
����a�3��^�
���U�ᘞ��+˘��h���G"�5��f;�h��"��s6��\r�$@�h
��	ϣ����A#Y�^QE^o����Bc+�7
����|lj?7P������rI��J��1*;`dń���+\6־8\�y�[G��X��,�l�Ao��O!���`>�����6o�푙�Iv҈gG��Q�1��i�dRb(��AilҖK��D�9��P�b����gU��A��F2Pn����#6��6G�B�8� Oא�;��zD@�%=s����I�D,�sLM70/�e�X�$�"+Q����Y=�0�a-?�+�0��ī��q^Tk
�dN`krĈ�=����r������13<'C�f$��10��^K�w^ V
���=nΘ)F���.f[[1�9�ƝmY��y�|řh��ܠ�	���{8e��^X��dt՚�x�J��h�.Fk*��j
ݩ"@���x�6�T#��Ē�n���.
c"U��r�.A@�������@c2�#@#�/i<�F�yU��pc��-��Cr�1
k������\�%�v���&�=��#�h]�jx^s1�I/UK"������N��W��c.��e@�9 5X'��2P//��ɀXbЮ֓=I->��AqQE�'��իG�⣂̧�2h����&����r��즙Y1X���(j	�"(��l�dCl�{ZG"�K�	H~+�H�ʦB��
Y�D��������r<��eh��6:8(�l��G���|OE4G*Z�뢥�X�B�#l ��h�	R��H�~i�dnR��ж��V�3�%�s
�h5��SLe��ĖA�u���S������A��?1w�e;����QrBC�U��P�ͽ>�M��t^��	XD��\jm�0�C���O�ǣq�mP)�l���"e�������/�,l�[@�w��[��/NS�4 	�>
۸u���Ƭ�:i�Ա����%��IҤU[�z8g�n짶Hz�Rk8,�̉�PC-�Q$�<�����F#Nb?��U�X�{���b�ʭ���"�Qè��+a!L3�>�шvz���4Y�$0�&�2�Yi�JA8�`L�Q^��`Иn4���c��˼b�Ǣ�xlя��v:4�������-[eJ��p��()�?�aV�G9��8v;��	�L�ٕIĞ^�����t|ظ6n�����&�3#~��{x �;{������b;��g<N̪ȃm9���t&R��&M��/ޥj�,��f�^�|g��.A��NG��^�W��"��QPs|�EC�Ӛ~��q0Wk�QUW�8�G��}Ypf+C��(�]�F�-gwU<�@Y���⎒��L�	<���(2�Qs��=�%hb��#t�J�͗�raA4r�UU�WmY*���2Cz$�`��N�}��jr� �p.��Z�X�����8�b�{�����"-���$�h��!��vY���g�� \��?��!�N�[��J��� �L=�Bŀ:p��Y��?�!N:��qAA���E^����YK;����h�m6�_{Z1�^��x �ZZ��6W�2n�bw$�(�X��RO��b�k�"U�Ĵ�@���2��j�mlajX�,(��|��.\��de���%�V�P�3���9-ǤQ���%�F]V�#s��+��$��0S�D��Ȇ����,Z�`h�%-i�V�e��nte��D��-��]&�LŒ�ԵK�=��@]�x�A\���fԛ��W��gd�]���_��p�E�;e��C䨠��` �;�VE\�,��~����@��ކ�:��@�SC������	Y���p��h�� %�!`�
�)E�i�x��³(�,F�h4@�M��G��b�*�R�T���a�̆y��)%	�k�.����}+SQT��)�I�+��"r�����aE(� �b�����Y���xW5�™,�-�}�E�GM������yn��p,�b`���2uG���W��r�����8~�B#��4���ҵ�g+�" ���S�x��A�!�Hu٣IA�h�*6EC��"Ҙ�H[	y�e��scW�cQ�����+�ȃb�?��NTXp��b�G7U�4�IHEJ㙂�x�ުB�����!zWd��"^����(�m퓖ss�V��v�5h��p�H�s<�X�P�8�VܒO.�R扆��}��v�s�X�	wR���,�#^���S-��E�D�]�㸳G�Q�jq99��yD/D�!�4*.���q	߉�J���>H�5��w�r��5��hFa�I,��,6����Q8�\���q�VBd��zRdU�x�$o+p��Oȭ6�xc��:L�h�Ck"�$�S���Ƹ�H;1�SӚ�]�,�f��)dؽW3�|e܁@e�\�(5Tb1[U��bYeq��xz�Z�X�`��!�������$��8�1x$0��դ�Bn�(pVK�\�x��ʻ.�'A��6�=��1���A���Z��x���Z u�:��w�`��f0i�p��5 �K0\�^�����9P}�P��-�;$�6��*v��OML$Z=�~W�c��g�f/aK!G![�@'���{-�	�P�6U��rn��e�B_�q��	j���y���P�3����(B���#1�#CS�C��e�X#�h�t���o\��>J9Z1Ĝ|@*�6�ۊ���-֥�����Eq}�u᫟�\;o#�~g���/��̣-F%#�*8bwt��҇?n�X]fkD�Ϝע�:X�9=����]�>T�9#�N��'�e6�����E�u)�U&��8Tۤ��^-p�-�a��Of��A���"�zMÓ���u��Q�4�џ��M[d�&��C��w��ϽL<��z�i�6��Gj^���1ƪ������%�F�g_��~!ww�Es�K�z'����-���i�]Pm�П����p�Tf�k0;��v��X���,1��-��>KZ���U�Yո`ʅ�X��銊�dK^���5[H[&&��>���_Ʌ���(�R:��}��m�g�]��x�����/GO�d��d�����~
ؾ��6�'��K_{�֩,f^�8���dԣ�j���[O�U/�/^�2�6�@D29�?x&�?�g?�J۩�2��^�y�Lm�Q����_�_��'��h�7 �4q˾%��Wc����jaO�
T�G��5l\�����$��8�A!gK3��M3�X��7����G\����Qk��n�����n�\�+)Vy��5�ח<�I�͙a϶
j��~��E3U#��̆vY�KC�h����2N
�KK���}䪲#1�2����U�`{b=w��k+�B��[� ���Ɠ�������2�F��%i���u�#IG�G���B{%7�S�SF���B%yr�ꮲl@ٖs4*U+$�5e�f����T}��j��e�㗭Ze\a�Q�߿ҋ��%�EVVÛ��f`!���ES��H��9Y�,;���^����=���.������o�#���^��X��_)����7Y��2u�NhT�L�z�/D�����Ci�<3�GPZ�����ל��u���MvT�n�����ǆ�ѝ�Ul�l�dM;�f:�sW�r���5 g���Z6.�U�f�#K��]��xմz�aC����Ov ��x�2f��X�i�/�հ鍜�}a�e�{�uZU^�Ҽ!ih�8��J�G����c��	�����۞�o��o�uzX�R���Fk��+n(0�pƑih{�=HU�+��`<��f�'�2��D��7�B��T�pe�h��,�dWOq�C[��zR�86��j3���� ϗ.zY����.>B4�qBϑGG��*6F��-X�6��\���3B�[Ȉ��s��pe+���ɱ_}G�T|qn)%��I�����-������Ɖ
�FQ�wN����윂�D���V�[�����١s�=_�ڞۄ�s�;�q'(:#V���?V�1֮[-Wb����2ʨZ���{��S�6%��O���y��-7��+��WV��<�Iן�5�IL���;78�����z��qn�iP��լ��<w6�� 'c-�k�v_OC3��3K#>aS���
˝T5���G��u^��aBV _�� ���|p�dJ�C��]c�T0�^�ޙ}s2�K�Ń��3�%�h[�}U�c#!M��B��%���᛺���6��u+�(�	'~V�U��:�*7���=6��;�jh�G��;\�N9�8�}���7��0���bh�Q���|��sN�K��h�u�����l%YTKX�HT���(mP�:��+��݊@�D,a�Yq��F�y�(5�9������w�E�(Z��X��aeO��S�XAUo��uP�;�2��Lk跢���-v�l��e��&4���U%�?Y����Di���r�Qq�,+��,D��!���(�4�oB�r��_�_N�Z~?�/�)U7�I8� ͦ������̿-�<�k�"�]�ܮrH�YK�c�M�����(�)���e�Ga�Y�G�]��I�`��W� ��}�}��4�c��љ�<�w%5�Cd��4�����u���5�m�w��ǳ�����}v�z;�[ Ѭ���q�A������w�,L7�ǐk-�Ά��X��_#��l�(�� ��2���Ώ������P+�+)F}DVMA�Z?����ֻ��*4��i�NT�-�����0���,/���|��~��ZB�G�ח��$'uKqƃL�I�-�rN��1��(��(1�n�[y�z*YD,��r��s~W��Qva�"��h�M�ǲ�w{,�>���Q&����O^��m`��ziM༇�S�*'WY��_23Fc�Mkڊo��U`F��ベ���a2V1Ũ�E;�wؔ��Ga��^�v�Fd�&IZÜO�<`�Yl�A�>&[���� �7����Jo�w��+>�[�N �w�&�<L��������`�s-��U��"i~��!����A.G��,!]Y��΋�}��w11Q�V,�.�(\s".�MD�-=���m��d��jv�{(�й��]t��}'&j��-1��Pv���sx��������!O�
:d#U���b^��ui2�]������%,����2L{U��b���N�aZI�f��o:�_N�������c��ba)JQ�aMI���LU��L6��}�6pE�>����T�0ꃳ*e�����KP��;�X�T�βD�<*a�4�=�������>&����W.�^�%[��ܡ�X�#�*b�,��M���Qf��>��Z�jb���F�{U��Rg��+��=:r�d̪��i�v���}�C���
��+Ǒq� [���̝�'
����U���51���`��2.)�[%���Z�2Y�`1+��P��x k7iCd���o��zݎvw3�Ċv&�<܏G��I�;-�W<�������pYH���1Zǆ+6�0��j�JcF����:D'�jMk+r�īh�^��(o��>ܰ%��z�ݥv������Z�����Im�ͱ�
.mj^����la��\���̚��H���Jh�~���
ƭ�c���G)�f3�1��%pY ��u%�WLElMd2���Z�]����N.�/�5�c�����B�b�l��zl�[��!q�f��'�Y����c��E5d�����HG�?ʞa����i��q?j�]E[x^���X_�f�z�5��|�++����ވ�Y���':�6F�6�[E��EI�(tP[��U�D�S�:�y��n1ºz��e�~��p��K+�L���fD?�J���,�8�N�;;�Z��5|
VY��&�J<�td�
dD���ŝ8��]폰�{���9>+�u��AY�V�W�� Ř���}z~����.0'%�sS5Z��Gꪎ�q��C-2He���E+Vo0ޥ�$�U1�3Pau��XSd+&���4�R��ͬ�5tF�.�b�Vv�6	��T�KSm�]��z\�'��h���h
�E���r�[\��v�-6�&������Mc>֠�Q��EaU�
o���g؊}&�}�7��M(��GG�E���{ޕ�-��mP����y��cj'EiN������a��I3$���@1��tǛ��D��(��'2�$����d�5��U��E�^֘fV��F(N�h0�`Ҩ?R�B��,�Б�Ԙ9ʴ���i��H�LB�S�90ΨA)l6g>�vߎUl�����(�x@D����x�q��H��^}�@��|h;�g��(�[-�T�`XYs��D�xP��U�6�ar���!�O<��� w�"�r4vY���uВ3�a��ݪ��X�����;�&�|�f�1�F�q�s�?�fg��.Y,O��X�^^�X-W��o!�~��J�ɝj�������"�(��v��������]���6��*e���H��]�j��)G
���h���:�*��l��#�0NZ�)n����qF}�"��^����C�*�o5��ׄ@xOfbh@,�O�4ǘm-p%y6Af��k����4L~c��d��Ǉ�K�s�����e]�0��m�L�c�*��c��ǸgF�r&��~��F%6W���^g��k���C��/G��/j�k�5���f�M��ڮ6�Ѱ�Q��B����jL�+rx��
i�Mi���Q�.�gv��|������k0����������Ñ�� s���Y�8@-D��i�X��*J<���:BWk�,k��S��f��G�w0]I13a�]�����Y��k����i[q޹�cv�F\�5���7@�kϾλ���۱Y�%�-Z�1-�G���Pm������hh�r��r��������bBN��x��L����Iy%��Yۨ�	�j��qе�Du�S0�D1ĭ�� RN�I2��3���(��.w�Ot�H%��Ii	�6M��W�;������x�_~����ٴ˱z�^��$���V|������֕"YS���	;/}8n;��-;��Qo�����8��4A�q�iC�D�f%,r�I|j��ʚ�0\�D�7J��v��s�@�F�4��¥;���M8`Ho4*�����KbC]�1�[-5�r1�'
UƑH[�p!�X�V��\s����ѻ��q՛��z�c�
䣞���Y?�0=;��z�x����o����}���O�7~�٧�;8�8m*�-�0�b�����oEy�c�T��Dl����}Ѯ#ͯ����.()���_~��#���O�R����@�*b-%?��Ǎoz�|K`7��JW���Ko�����0�˞�r,UN�(n:��,76�a�y �A(F�ᥡxm�%$�Z����8��}�U��]��k?��wnr���թ��:��=d`�������?�?�����Y��F�L,�50Ԟ��:��&a!������]/8\��ڒb��a|卯uu �6;�|n�1�����bg��KQ�r��-2�H�bB1��kk��,��+������`�\����L�A#Ws�+���D����ȣ~�"saU'��v��tw��O��M�۵ �#���,�1�%�R�0�Z�T0מF֛�L��x��G���6b\=� �c_�_f����8d�����W��w��k��U���/�����Tis�ץ+�TE���@0��s�ծNe왠$���&�Ɓ�:W�}�ӱ{Ǵ�0^D,,.��`��  �:�����u�=ޅ����	��,.��,?|N4����:K'�@!������p��	`dq1���dQt��+�VbɤV�"di��S�aK�ŗ?��x؏?��P!&Vl�),�D�q���B �@ql%��ۿ�CK	���7��]��,|/]W
�}0ֆjE)��������T�Dh5�sS���X�$Y��j�1e�]mn���-.��"���K���˰�T�⚆À� �z�D�S�������+�6���d��,ʩB �F���gl�o������ܪE���Q��~�z-���(&>���!	[M�6y����|�3��~�|�s��O�|/GufZ\�B��x��d"��`y����3���R(�>;�"��W,]$.8��LOOc~~KKK�29<6�Ɏ����D+�Sf;�V��/N s���U��"@�{�^9ƕ��*!�}���1ը���V���w��� 65]<�I5lV�bJ@���G�����Ǩ�V:Ǐ~�ݯ�E>�=�hO��ngQ+��j� u��V����	-�c�!����E*\Wq&4�Yg��Zd0�(���f�]���녣�U����r�\�;vh�Dwq���H�$n,�6���w�]�y�'#ɓc^��lLo����Gr�d�{�5x�c?������Kt��0(�������2~����J��Z͚�W�B1b����ݟ�'<����A��ʱب��*�m�~���qz�y
��%��Y�R����"�B,Sn�ZՐ�Xҹ�D]aR���͊��:�_cȍ�s��W��5>�G�+b�h�'�Q�gq������v��!� ��?"�LLg�~�C��O�5Hn�F4G�i#A>��X��s�A�f�������H�!���~�9x�[���={6�G��2��r�I,��]�ڡ�J�ȴ�g?�Y\��������fu�J!��ح2<��T;��q8��v� �4;3��
9 �L���©��&�����׆;7��׾r�^0���Ƨ��SM|e��(B��G~����\��wź�UMQ9�,��	��6Ÿ��E%GV��U(	��2ţ(�;wlBk�6��zl��n�� �S�����ᅿv\�(Z�%Gk�`��H��SSSG���V��^A��v�: �D�)=��� ���X6��Wr��䓟���k~w��\Th�E����Ck'�# }'ល��O�9S�����¡��е9NqL��ۉ�:���P9�+2*�+����_w��fkZ���x��Ql��b��9���}Pkl��%ફ�£x>�h�ǜMX~F���dn�U:-��^�?��G�B��)_S�щ��s����6X�B +z���y�,;�e	����O�����Xs�ꈰ4KW��qѹ���������%Í\� 1�Xͭu�.X�W��TN���@�	�C�4��G��hvW.�ԯ'FZET�pi �0v��c�_Lj�ȴ����~R��s�?|�׷	�]Y�����]�� ���I?j�8��5�4�fx!e%:��k�������>|<��'�����Õ�������*w��U����"Sm��Ts"��ߍϊP��L4|	��y0��6$*�&]Y�ǔ��=�d8�,C�h8���0N�/��ึ������K��+~�yY��cbpM�h-���ʮ�m��4���F��6+��:�����E[�k���J����1�!(W}]N�Ĵ�ߗ='r��a��@<��n�y6�]8&te�_�n}�(ߺg��-�5�����(��&�U-VV�z�&F{����J��v0��J�ܠ�*�ipj��q�rj�D�+
l��D����PR�zlGDLۂ~�ų�AO�\���Z���+_�v����U�A�3ϣ�+�׌�`��>�[vs%�!�[u�z��~������7��O�w�d��/���<���1�Q����W��f�b��.yG���u7`���jk���MOa�)Ζ&B�+yI�ڥ��k�7y�H"~O���q�Rڷ>C�B�;f��M����;��ٳA�c�Z�i�8Q��]GW�b���v]s�r�s�N÷��C�lQa�hvO�=i��U����%��佒��~����C�B����u���B"5oU/a�ؤ:@�Gx|�T큲L8X������_�7�.����遟�.�r��VL���V���Gj�uUz�
����V^�q�E[��I��k&�F	enS3�J�=����Z�kaLIf��W�����˗���<�"-qb������i�b260�7��e�T�r������k�ť�x(~'ݭ���G���K� ��?V��e�	Q���G#wK�1M4D��9����'��߷�B��/����ԅ�vaf�z��Ny�6��5�e��� �#rC�;���P�� 8v�C&<6nj^�a����q�RBS�#�P��Ʊv���Yl����/��.��C�-�}��a	rd�� %�*�rKN�
�:T���	��S���uo}����@�ܢF0��T�r��T�
7���Ϗ�j]t�3�D3�L��4�n5,?prV���=�N�3�\�	L��iL�X���`���5�̯}�B���i�a��(߻�?~���_���k��!q��(M��f�{Y>ծ��ط <�g��e1ІU_�k|%�Kp)J`�������4��zJ�{����	���7���"�G̘D5�S���D�&=Z�a�QK�ԕ�e��!��߲��������[���������]�e�Y�%-f��n�[��;$첋��Bޗd�v��T&���/�G�����d�ғN��=뻡l�R�"��|��/�%�_��(ƅ���:��`Y��XV��h���k5,f�i�$.�]q�Ȕ~���.6o9�����َ>�����=��.6������o�lR��_��P��U*H}dB�v��`�ⓞ�Bl}�Oc�3ppd�ܲ�D���(���D�f6nV���?Q�梫��̳X�!3�r<uʌ�
�̕GM,�����S99�yX�s ���.���������蒋A����L �/ڍ��QhB���EW��NV�yB�=�]NF�2�����T��E�lۿ����E����^�
��߾NT�����5厐P�C�^�2�z�"�*����"�k�	��?~����#��Jt��R[�PQU�м���G��J�<�����\��G/:y�*K	�(���,�3�0�w��OL��o�t�����b|�w��=J�F��4����"p@��2� d�l�$V	eg���S�5Е�Ui:ɚX�����¹|&(j��/gI��P� �Bԧ6���,pѣ�����7_������YNR�{hb�c1,k>#��g�Q��[�x՛ޅ���7�G��=�OCM�)�$�C�Pu��G��k�,��KAT-X3�P�@�GvnnN4ƒv���ڼĎi /�]�6
ׂ��\�(C�c��p?���v����+��
�R,�Z-h�hX�j-��<`����$b"PRa� �I�"Z�0S�bkD0Y�^���/�S|�u���7_���b�T!b�E��}>4�j��V�/�O^�B�����|����H��1�V����u�@���ص��%䑙"&W��sG:�l�����w{%��6�T�v�T�5V�?����S���:�#��*�\w��!;���Fy�l�CY�Ly���RO�>1���� �Zؤ���#�Fz4�!Y1��.ϡ�
Nc�1:�Q��Hda�"�ڎ��<�E������az7��m��������z��
�ۋ����%������`�9x�o���v��IQ��E"�X�A�K�lP���!�C8��*��`Q!�蛲��Fg]�����P���nʤ��\��{�Ur������Z��f�20��&� ϱ�aB;첱<)�	�յ�-TV�*'k�7.u�|F�?��~���)=;ϊ)<���ɉ�]��F0�"�T��dd�!�HH΅��`���~?�x�q6�x�ȿ�7�x6�����`�i�7ƕZQ,�o]{>��k�;��
8l��p�C�{S{5Y���w_c8�g%܂�Q�Z���"涊��xdvI���'ی�,q���B&�R�,,P�ƐH�]�j!�Ո(�#��ȵ8�e`l6��']��+��8�.�RXUKк�X�ьR���Ri�j��-�"gdC�}�mŰ����k탇(�G�4S�E�eYZ�f����[ο[K��;o����x�k� 3*������Q��坿o����z��6Av�p㐣�	�F�11���L�3�9��xt�8��!c4g��8A\ Q@Y�fiZ��n���������<��}�{o�UTwu���)�����}��>�������Y�S6�$��'7?�=[�Q��n<��@�V���[�K�#:�����X�.:��U��W��V��Z3]y�����r�)1L�}��F�y�ݻ��k���UW����/)x��d�u%�-�j2�8�/�����m|��FB�C��O���9'r+�Я��gj�;�뱃���	����b�1�������/����1�-��Y��Q���*�l<��߉���S����ִ�҅�ƙo�0���7/�Щf�hh�X�s� �tUL=�#D�n��C�
9@SعR�8eۖ�"�g+�
n����_Q��9����&6]'A�-i`�QIٜ�1�K VYr���L�1m�&Y����O�"�%Gp��,�
���|�T��b�`"<���B1�y��@|!�V��vӱ-����V򒁉 koK�MOs1e2�`GC����K��d�S-R���S�qj����s_KۏW���r��Z��o�a/6�� �<wi~'��71����<�M"��
�JϤ-=�>#�v׫"m�X���|7#Y N���,�(�\-}n���	�DcV�R�`�Lf-�r>5��٘E�O�3SYe�FE[�C~r`���,�?�h�\�˼2�fc��v�1e��z��(J�J�kk�P,Y~�,���
�;��{�4)��/�5��cU�2����b��yM�Z�G�{���C�X�Q7%�.������l��-C�kj�=�^�L-h�-�b�pS��4NҾ5���e^��⏃���1m�8�������tn�
�1�.?,(>�5�S�ȹ_�M`��g;yߴ������b����l
�1Q�߬%cA�e�kMy�Ai�vD&�cx�J��-Y�mtd�X"I�E���x9C���&Β�OC�g��
Lr�q��5�{�հ� bh~	5b�,����H����	Ѧ���b%�ܻm9_O���!d��@��Bƒ�J�f69Y��U�4�
�K$Mc�6-�+��s�֢�U��6���t}�7ѥ�S^�d�X�}�z�6`�َ�	L5yv������\�/;�b����-up��r3������	�Y���B*JS������#!MS?��%�Li:����3iS��&Qm�jV���B�3�vC��3JF�A�p�k�.���h�c�v�L�u��%�,�����T��!&@�31O�l;��a�)�.�>ĝ�:jrjU7��e�l���� 7���+��a���o�
8�*��9G�A�RR�����rt'J{���MN�5��d�#6�ݜ��\a�d�D,�oX��;&I���3g���|>Y ����b�R�W�ТN���|[A�V
d��V�Հ[�+���u�Z2�Cc��:-(�؆�^j�����P3ju7;��6�u��!�ԄWC3a7A���0y�s��	U�0�N2�EExZ�s�����v�VdbҮuqX�{E�|�oh ��CՕp�	&5Q�X��e�f~��U'��z���`
����C�,��g:� �5���{�&��Ս�5��&,bm�h��h%�*)lH߰r��]���\�G��y�ͭ.�\��:�x*�sZO��vsm�@�+j���� �3ϓ�|8�Ψ�E=Nlu��mi��,�ew�|Q����r�)�A�W���%	��+'���k�Y1���]��
=�]�MPP�2�'���H�$���Eiw�Ԃ>hT3	�e7Α]X~f"�f��R
;���H�K^`��.��EK�ƒo��d�99*f��
�Ŭd����&���S-~f��XJ��)�f���Z(����y�٘yNgi��&��{�\ܥ�%	'��_|����ر��^)h;�o�P ITS"�Q��Nd�+MA�X$���b�,xWI��]C&� ����6�����{p��g��֨��/U�5�s���3�����q�a �-v�)}c��5_S;#*�}^4aQi��鉐6Zu�Dk����h���B��<�>��M��T���+rltŪ1����QI@�YO�H�S�/yH�eX�wԖgU$�<��;������d־�\��W�c�J�N�&bKw#���^8�5XV��yY��� �cS��P.�B4B�1d�\�2�RK��I��GP7Mz;�#���G���xg��4���Y*:&�T�B��&})���,'�MY�xj�b����x�ٽ���T��^�Xhf��d磂h���aW��]��y�0��F�#��"�%����a��5Q�IꚲG򋤖��H�%	wD�1������W��b�T[y_"��Si��B���٢���!C��G�g���*ʎ���F�HSi�S���MZ>(����ڬ&_�\6�c֓�4�'GFsF�rX^'�$bW[����N�7�7}�أ�:T.�Y�5	.)��/��7ɸ/bkfy��!,V"ylcnF����kI��`;09n�r�����,(�ʂ��y4��-WV��/��r�䰜"ir`����,�.��9&�����Z_�h2L�6z�&�`��;��P����U1�`��VPk����#aH!''psr�+^ ���9���rbB7gw��U��;6�QW��ب��j��ۗy!CEu�T�33"�r֋�*��k��&����햇ju\ k���1�����/�!y��'�]��T�sZ]y���VQ��\��}�w=fL�[az9Vrh�Mc�%��ИhCu����(:��%���"��u?0AE�x&�M��=���:�
9N�{p��c8�����0|�i���-���<�\l}�)1	c�h�݁sљز�Q�|�|P	�e2j��a��2���� ���5�#��k
�a{W0E�1"��W���k�И�����ĝ�������Gy[f"�ΎB�w�F����ry�蔕(��("X�>���{��`���t��L�,)�;1ʲ�W!��Ƿ�<6!�{��?N<q��.��8�����W����/���-pE �����q�Y���'�C�<���"L�\ds8�2R?Y��XL]����"���)z=�eQ����L�8��g��W����gw��t
.�����(�[������_(��)yE=���k���k��O\��\v��j���D��t��Gb�Ƚ�2��;d�����k�;	����������F���������^�w��7��~��r�;X7���{���{p�+���W��ct����+�a�N��f�&Wk3�~�p��+RS�없Dc4�r���~u�����K��{o�[�r%���3����%B��޻Lͅ��!���YGs��5o&��o
�'��ʳOö;͙��a	#u��h�Q&�TZѶ��M�1ˡkhG�J�d��1���P|����ӂ��������o_{>���?Fm�p�ӣ�n�S!�>4����?˱*��=�c�����m?��-�&&�+�1�u~م�}Er��D[��;�߀��0���"�I�"��B��.������L�;��s��-�:�����!f��{�O�Dy���ˏ�	�굸�~w�8(J�!|����g&����v\��w���l�	ڙ¥g��~�;�\p��w��ߠ��l��s��1��k~�
����}��(.��;V1G���.$QgqGփ`��M�D��y�u�Ȅ5j5��qf�8|j��ȏ��^DZO<��%��wn����>Q��h$f��\��	/74�6[CT}�+���(&6���^3��*:/Ml+q�����σ(����+O��:'���~��9�:���ߎO|�2|��7�L5߸ �07ׄ@̱6u|��:�k�|�F\��Y�M}b�E�g���$��Π$�xσ��o��ٯ�ת�������w���;n=�Qǋ(�R4���U��tF'��\���rΠ�Bn�Q��:/�����]w����β���׏�=덣�W�O㸕�䬔�#��[�S<���8���_�"�H���-y�zm�6[*!����ΐ�jc�R0)�ֵ�v�Gan���D_�,�˱t��S��xIP�`���q�
�:���߉�U���Wn�����������D�4�z�E�4��T�ڢ��N�Pm�ͅI0I�&���#|5<�Z�Q����������.y5zH �h��a`�����ȕjJ�ҳYKIN�Ǟކ�_�U���7q�2fĢ��E^/i8N|�\���,����<�� ���y6�����j;vlǘ�m�=M4��q�ƺNǴ!�ã&�W^7gń��l����<*��J�*�OU�擺Y�p���73!]��O`V���Ę�B�%���7ނ�Gc���R�c����0Z^�����߻_���`ƟϠ]$O$�Q�+�=L�މ�+����4�W�*���FPA^ݖuuOn�!��\��a�9����w��:��ΚXh���v����ג�[y�Xe9L���E`b:��RQcIGb,�%Nn=��X���[(���"�ڻ�ֹ8�k�u�n��|5pꩯŽ��BvbGk'�]�m[6c�3L��p��ER��KLy��Zr���u�8�4tF?���X�UJ����b�ú��bӶ]芠޽���J���VKZ%����v��ǛE��
8&&�"���|^�g�h�����q�[~�ݹ˦��"u�%=6@��v~35������;��4�7=���j5yt��wc�Np�l-��gZTc���o^��7�{����X�Z0�Zq�H�\��xP_�Xr�Ĵ��m�,��a�7%�r<&f�f��L�?�p���l3�Yg�ؽ��!^�oz��}'`�ګ�G,�+.��>�"�>|9N���e�0GrX�k�i����Z�ZH��t�n	���؃�}�
��0�v�Jƕ>�NΥ�	f�9Y����u_��?��I&�g9�¹��A]>�����o�����;Q�2b�#u�G�֘�1+G�H\�T��b~7�|>��_·nK46N
��]�㲋�����n��j/��W��y�w��O\���x+yR4�tξw��\���%\�\�Șah
�֓��6BKH�J�,z�����|6?��y��V��A�����<��^��?݅��;kN�㺯��]�?
�z�L�|� �;�߅�b�TG&ЊM!�U��N
�ɍd�c|r~p�#��&�]y�&��]�ɗ��^�-�o����L 	J(M��O}�Q�Ys<vEں{�z�$������	<��^�i��V�1���em��h��h����Mw��-<���P[G�-�?���pʩ'�7 ��~��=�1���?�c�uڙ8���`/1oxRۓ�z~+J�1,�^X�8�Y)_�c�0�����J�7[������U�}���Ҡ
�6nA�H�}�I��ûerD]�{<Y�T&��z�V�{�"Z"��<}�����N�yL2-�X�t#Gf����t�FmǊC��ZA��06=�F�m���y��&�{�!�6b�����>�r�iN4LՕ'
0���P��N/��61���c��0��Ąn������ڔ7j��ʽtEM<�m/���S�L!V�	�� (O`J��]?} w���L;�ȊI89G�[���s�a�B�n��b���J=�.*�5��07�f�&�Lݣ�95I������SutR��YdS��Y���4�b�QlZy���8x�X]�ZH�E����f�V��� M�_!3�=�Ֆ�ntM9�b`�R����{O���k�e�6�aƕ��[BI*5yF�¸��W�8��mkg$Zn�$���wCK��_�Gb�n�BQ*�I6�6�r~(����n�����8>����2Bȸ���TC�j�m���fՙ,�/�P�%��[��$Yu_A$���j��9e5z��:���lƒ��<p0�O�g���fFj}v�����hn�>r�os:L�j ,�,#�VEw~���S7�8��s1XRijK�L��.��[(��+�6���8�9I��+Ô�P����@��*�дgBNfڇ�R*[�]	�ѫ+IM	�YN��k�H̸dȘD��A�f�w`��v;�?D&}/���6|�,1]1m+%��wuA�W��>��,:� �.�9r%���P��"*xn�/0ĲH�%�i����3YעB���1�"_Y/X�i-ñ���Nb�gW+�px4:ME:i��r�C�%�]�ˑR�g����4-k�|6���AH�� MFnv����L'1�_o5ܒ�0^��q�E�1̙��>����%�D X�����m,??���n�G1/��4�5��}�}���[��(�=���0��~ـ����I�Ք:h�<jXGܙ��_�N��=�S=6`cv�y>���{�s�[�����g�M���Y�L�C���Z�GuxT3��-:bAl�n4�I�T��w�ƈzi�� 2ZG�3FA�^]�����_Y#k_���Y��K��Bh�E%�d�%˲���~��k����U�@�ڲh�bT��G2�)CLb;�?��ɩŶ�,�~i<3V���|��	5�[�N��~��:�X <2��,\ʉ�x2��vD>�P�F<��M��^̳F��l�'X�7�XԀ�G��K��YMg��؆S3�dwT�t���|�������}��2{� ��^��J�wy�PALu&�v�Y��ǒ��,�a�t��J�����f�h��ҋ�9�\D3��i󖬒l@�M�`
۪UK����/�ݬ�Yi��l�T�~��lz��m:T�k5�,�\�[�[�i�X�	��y�ġD��L_��L&��TL��M��fǓ&A��ep=��\7�f��$j7�a�Sd�Q�PP�D$$E�m���C����󥏃���1�ť���c֏r"S�?���5�f[i�>;0˫c��E���O��n�8����3� K��h�2��Dq����[�J3h��.8Øb߮:�l����P��hE[�0Ɏ��T���5�A0�\�J~_Mc3����J*3�=����Ũ�v���Psj�\�T�Y'jj��tvvZ��e�Y�+�0$p��.c,�����݁ߘ���R�BFJ�M�S��I-m�vc��u��j�|l�8��i�]*U�7baP�n�,VÑ]W�(��:äh�h'�����I\[39�HLN��&GՋ\<ϵ)�L��h���	]�^�B�ߑ���g����#U$Z����=�1C��Sj�����g�7�I=F/����� s5us�����"�֎��쎒PkRY�C"�?��ۊ�]m�j&��x��<�Y�K�+:U���k�t��f�f��,C��5���c�%L�%���Tr�^ʤ�G'He����v��R{�� c#Qqj��z��w��ۨ�b�G�I7����`�E��8�'aI(�t�~�i����1��uy�jf�.���jO[f�����D�܍Z�wш�9����~Cch�]��fn�5�Pt�&�DU{����/�FzS�jo_�s�xz��tP��Ư�g�!���j��p��?�-O>e�J���e�%�ݘ�1��4�3�d���Z��\DzL2�~���$��a�Y\��s�n|�~�j�l��Ŗ���0��B�%�ϬtP�{te�eT^�bM(ܱS�����SN�\'���$J�1l+δۄ��4=]t���B��	�X�UC,&��f{�+VL`�ʕ(TC%Jcy`�e"������ڂ9���V�1��;�Be���W��>
f���n��L�g�Zt�E�C�d��I�Z�Ƥ��zH��q��VKwp�
�U{f"�l�TK��0u{�ڤ�1j��hʢT��-|25nd-�)��U��wH��1?0�5��G�O�n��<׀�N�!ɉ��P��R!w�[�$�J���!��APNv����Z�S��	v*��FC�ZM�����[��<l�!A�K#�9,<��A�M�7Z���o��p�f�W�>��
Z�϶��rrg ��)=�CH��}�J�{B��s��'iڗM�jm>�(�M��e掺I���	��YE���ؚ٬՞�<K|;}W׿�wA�"��Ts�m�=ǦO:�ݲ���B�S��jwǦ⩊�S� �-��p,ڎ`�PS���L*;�\Em}v,�r����N��_�l�Z� �g������ɤ�ϜI�`�g�zb,&�Ȗ���v���G2�ˬ�h@S��3<���1�*Y2S�Q�iE΀X��Ƭ�����hu{~�Á2<o!�J�@��]���=�6�<ƞɈlNbx*L�(GU)���Sx�hV��v_���a�}��n���ps�0K%����K�kL>�)2��*�%bIP�źP>V���׷�%��d�Y}��\���U.>���YI���j5EӸ�T�U�`9fU~��'8i��4ѡ5e��quc��D���$Y�Q��f����4�~^F=f�˘m� ��1�	���`Ǟ��9L�U�]M��,SW�)m`�bH�*�}z��2�s�d8����KQ|��U��٨��R�\*��@�VIg�"���)���xP&Z�`�I�Q�X޳���S�@��ݘ�������A��C�=�m:��i�����g]�f$ڔt�8gI�.�(a�gԣht���he(��j
z��,S����������ʨ'��MicS�d"Q���A1fيI�P��pkʱY��H�-dHk"�Qά���f�i�bF{e�:�b�ٽ����1��Z���O~.��mHfg�b��"[7c�.R4t�PvB�S���gFN,���4��FMP&�K
��{��4r�u��{�9�t�qfy}qT�gO�56|����~g>�g�����=���
��bQn�>�@�'�t�5�fo6��o�Y�)�\s�k�m�d ��G��f )`B���S���ȏ
���=�B��i��a"�@�0--w)IV�jg��0��3-4Km�je=B���d^[	Oש�B�u�NS�V��
Y]�$0�����ޖ����2�$0:r#�Ly��b�fy���p�H�e=�M��3t�Y� �D6Dq��
�m�HyRR�Fj�����ܘV�i�΁����P�ˏ��t�m	�����)���!i�l9H��OTS�-�Z����I���+5�:cΣ�.Q�����NK&�.�2��_��+�{�pjd��[��\�<fe#EE>��06���רFI��@vl��x~>�D }8�y>'���b�_������J_�fTE ���$,������Q]�mnik�x5�g�@ǩjL�����S�F�l�+j�԰�e~�����*�[Q���\D�*������{�pN�4�:ن<��X��.�U��@,'1��b�9%�˫А��jH�|�Y�c���g��� G��`��t3�4_�$�4�i�D3M�}%�=��E�@D�1fs�����	ztݢ��rSC���RfB�D d��_�
x�����j�tt�o��;��m,]o>6�GY����x,�NytT�挋5|m���pJU�Ϻ�cȻ��E�p�Eb%lD�Qv�f;%��2�8�o)��9���N�xEF6Mb:�XFY�܀����9;���Q��M8$J���&|��;�"��l�*�\���Z~�d��d�A���1�;����_�����j]�p.��e,'����Q��I�I���D)[)�4/�-:2�,��r�Y"V���7,s"�*�zu���� 8���u%{N�k�
�d��'M�O��f&����۠)Hb�VB�9�T�ihW�*h�A�(���ޥ֘�?���$�+0�6!/!���`w欦�65�ɓ�yyͼɵ�^(�/C*|Ij2�� d���u���NL��TK�r��Ӂl$�.�3���0f�%�R�JD�%���s0&���G`�,��؀%�z&3o#G�5�-�:(��+g��/+/k/�'�0ǡ(�f^�C����k�(w=8��7�'��Kר��-��p�Zu+k��t"s�U��O�AG@n>ߑ�5���"��vC��	��0A&(1�SqR�������f��O6�Y�T�+�u���ԛ@�SG�K����䞺ih�H�^W⩮�0W혓�(X�A���`�.8�RDCE6M�`�]�-^�G�rd:6�L�w�ɵ檓�I2_ej�2�s�r�5��h�S+�y*0C��ɤ���b��b��Uu�%a����[�=E�u�[�9����u c8j���cCs4���|�/��#�8$d�]4SB����=�;m�}B�{�N�i�`�+���Hh8��	4��8�<�иè�e�ш-���X7��	-'�̙�Yģ�ڋͳK��Ԉ�蘒��`Q�}���ibx�X	mG1	���E^o���3�Q�T:�}��"['��,�����Q�nhh��:�M�I@�fV�(��\��ȘoZ��(�{��q]ߓ#�����6�v����5�FNO(H����b���z"���Wa$ECО��B�]��X)��2�<�ג�9����O3�f7҉ɸS=]k"g�+M���?��S��(3a$Z����d�b����	f{�q'	�'uc�IO��H9@�U���J��.`d	�����O�V&b1@�s�`tc�\7�ϹCb�9i�T�Փ�CS�x�ߡh��Wn^�"Q��y?�Ė/jy�Q��p�-TGdG5v��D���f�i�b�;���9Vx�DF!���5NJDǸߍ��|�:��sI.g�.�0B��F��]Y�Ey�1�gŁ��j<�q��0����h��>�h̲mu�K�����{�%��A�a��e��1���T�݊�ĵj��YBN{'	،v� 	��ߗ�):�޿c��C���׼t^��r<G= ����~�|�=��m�[��"�yG�۠�.�Fԏga �!���W=��:k��� ��Ҵi�E�p.�̟x�BŐ��ۋ�ʊ������H� I㚝h�b#�^'�B��=O��@OuQҸ�=H��5�����������S�v����Ǣt
�>Wұ�fKE��g�G=���C��Tk0�<���v|�ǳ�Ug|��z�0�[q���\vT>�|Of�4~��|+V3��h1�Ӗ�Ԛ����
�o�ƻ7�MC�9\ks3N�&?��������a�El�LD����az�?�隴��/��;�FF�l6���O����?�p]o�k;w<�X�Vav��7O�����-��M���շ�cc��x�ٍ#pm���6�s�|�������_L��%�\	�\��_�η�������������߽`>Ƶ���^��7,w�,������۱�T������9�\p�,�а��r���߿�'����ј]h+���^�����6��f�v}����N��/�(�l�Y�c9��P�0�(��8��_��:Ђ�a�S]�k�A9�ꄫ
��rX��2/?����A��D�B�GqS����Ǳ��)�1Q��e�x��I	,B�l�Q����c�ޘ(V�rf7��/F6��wʬ���֬Amz�����n{E��n�y��W�57s<�q�K�D�^�Hշ��q�qL	F�T^YL;�3�U2����ɏ_��|w(_*�_��bg�b�8�4ʗ
y��d�/�(�cJ0:����8��b���0q\vC�>�sD�'�v$ʣ�>����e{�cJ0d��O��xK'�\�p�z��ue�JQ��'ը��7��q�	�<��4M�M0r�eJ���/����a��A��˭��֣z�k�����Gl$��KO�^�؟�`���8�#]47�aG{.�0KGq�ɘ7D�� ?�C�����R1����O?�`��w�r.�����V����hjO�G���ڗ��Xf�8��_�c �l� ;vY����L	�Qǔ`�_i����r^�c�1��U20����5�����܂1o-^��c�s}�Dq/}$Ird,|��_��1O0�Y��s]�h/����e�d`̋O,��V�����Q�,�bj�Ʋ�ǔ`d~Vl��5�?D�Aļ&��I��|�M������Q���.'���(��m3�	�V����jy�Ϝ#��.�qL	F�[fa��o��,H��lCCCڈ��l.[ȟ�����5���pS�Q(��Z�P4E�NҞ庶��z��Uv�zY��-��2��cC�,��]�V��Qǔ`\|�ş���V��eq��1{�r]���/���۷�#BY��7��n,���K�X���T�3r�8���6�o����q�eU���8Jc�ڵO�ǔ`d�h��c��W���3j�    IEND�B`�PK   ,��X5��<O  g  /   images/c0642b64-198f-4d8a-96f5-22ba47d3499f.png�x	8�m��P!B�a�0ƾck�l��Nf�1ƈ��O����:�}�,3���'"#K��NQ�o=�|��������������w�׹]�u�w2�ڌ�[��D�-��8��ᄧxh�0��	��H�ۙ�Q�do���Lup�9� �������S�@)5���MwT�]�(vdD�?�\�	��]��u��K[���mT�
+G�yK}��*��~,�[��>�_�5��R��-]�[�Gգ�/Q�y���_��{>6�;g^bɾU�J���P���H��d+��Vfɮi�JÌ�x�>�?�UPUo*!>'�Y;]ʓt�m�ġ3�-b㺔�Ur��c���sX���^ς�cR	�'�&�q��M����_M�m�<`�S�|g�?N���	�V�{l�Z}.,���t�*�O��8���!;����EyZ��w�	")�~x|83纀ǵw����摧+�9˛
�h)Gbf4�'�I�Z3�����/r[C��k�.-��~�����2p�d��43����G~�x~r-:�@�󧨏�	�P��EY7⅟�'��65Z��ت~wj��C�bS�Jiw�0�I7R��n�}�Z}R"��Q������pT�^N�aBX��l_t�FD]Ь�#���v�c7�����w	`�r������q�
U	Jq��-*>�Do	^w�uk��[�^��{�U'�M�?/R#��J��[�bŅ�^�1�Z�G��w�Q5_�~N���g��~�F;�1x��䌞����jv�9&#:u�Գ�j��*���;�o�qk���^}����-}�P�#��o��f���)|�-���X������gs~�A�b$�I���[/�_H,�[���o��~k�����Y�ϴ2kφ�7�C֩�ʕ���:�&��c?ښ^GwD���nuc��ۙ7��^)@*Ƚm�wY�u,R$�`=�S&���i?aI�����m=T���qy���Y5�)R �GH�yIM�l�nVrdKެf_��rp@
�q\l��l$xY���M��C��ې�);�~{]{���>#����*�}�D����k4���-����p�Eo���}M��l�Ǥ҃_Y^�Od�\��̏�\]�Qm��(��n�{�l�8��4q��y8���;8G�h/'0k�[%�����[�[k�P��������hMK7�el���7ܮ �Sc٨Q=��.ubo�I� �Gp�fe������g+K����%{��H��K� ,�Ë���=qx�?2��������U�	��dD �>��A���B��zap@ 	G� ������a�O�p�}���B(D�h�v�B�O�q`-%����2XKG�S�[����VUVU����T4��*pU������z�퐦�fz�� ��BCC�BՔȁx����LY��
Рp�G�?H��$.�+�@!���;}Or0��K!x��\��_�|���T��a���0�����¿G�y���7. 8��IX/�G��S� ���� 2��C�oD���WM����.$��� �I�?����8�.��3	Ԕ��w�?A&₂ W# *������ 6/s
.@P<(?!�� 6�@�/��q;3����	���7�Q�0��3� �築T������,m���'q��2�+�jPU5��\C�����WV�jE����-T���OP������z��Ɂ$������!�8ΏLHQ�G�9�����# �� �S++�����g�D@ ������izzji�@�pZZPuu�T�ӄj�p���**j��G���w���x��p<?��x��������N�(���_K�w�כ�35�^eI�G�E$����k|���?��/Xٛ��3�6�.q�����)���Yyx�w(��������
�� s`�e�_���K��M��O��t�.�8@t P���Z���̑F�0��<�$��C/e�I������q���H`J9]vYX�r�b'��{v�]A�F�$K���vr���1��<@��loM?��@�����������⑻�6_lq}#�>Z�9�ݴ��`�V	N�Ɉ�O��G5m~it��!�H���mL\

y�F�5bmE�~l�q*%m���ɤ���y��+�Z7�Lo��:�8X�5���E�rA_1��ML�[�u���9��o����¶�Qff�);���=�F�u����t��.��2L9�����G��=>}}+B�aqt�}	�6���7�b����g����Gغ�O3���7C�嶷���WҮnWK�Q�a�_�EO��.�o�i�&V�b���617�=}�������fi��u�{��o�,���0�{������(?	_}��ڻ��E6��v`�����������?�WV�����l�i�؆�>���+�-���{u�%�)���PuJ�$w;"�#�2�S8��������(�Z�@L�.8o�����o�*����ϯ�'�\@����{=Ș8ܷ��7��-�%��+����e8N�=rfZm���X9�uƥd*	��5���g���r��A�?��~l��$x�w��}&�����6��>W�zw��C,W�-TTWy��v92cw��;d����h����`�l����.x�J�)�ą���{e��(�H�MO����[��� �����99:�[���Gx�x,�y������ثu<2u#ꢧ�ԏu �I�\���|�&6&�&����ۧϿ{ZY��.�װ2��#�ĩ�Ds[y�6#�UO�G�v�t����{�y�h�BM*[W/�R(�x �p��K�w�
�h��Qh{{M��ZX6���]W+>W�s�[Y��5�	F�Nf?֜!���vk��F�_�̬��j��gU����
�Ǉ%+<<��EQ�i�M��b6>�L���zf�J-�����.#�j�_�ē��j�H��cIl´��d��Ne�H
��0�n-�������p��8Ց�!�E�WK��Ns�Wg�X�����DҔPHh���Ř7�l�2��`�L�K�L֍�2ѝ"�5t��6�X��(w��c��{���]B:$sY,OU�j�]^���3y��8��:Qa�&f��7�3ya��
ZV��t��I�aw�,������C/"Jrh$O��i-�M�[ �sZ����;�%rt^ߢ/g�hȯ��P����1h�#*RI���h��n�Eq�mE�]���q� �p�-:���i��ET�5�}��2��r�:��COm"���v����'-��4���yQ1���JR�a�!�L.�sֽ�/Q�%:�6����X���5�|M�J�c��8����J�W�+9�^ɹ�B�-���h�H���HΥ�����y�K4�)SR����OR2�G�:�H��W��)�={֓v�2y!.���b�s�Z���������jz�BVإi_�)"�`h[�^�]�ɮG��Lh���4nꚞ@�'I�Y���Ǵ�w���<���r�#���󹤆&�(�L.�vE ��1�H�k��#04��_���z�dJv?B��j��%�{�����8��v78���⨮fm2m5����<����s<;��l!so�`�\`���K�Nz�q�f<I��	���[Q�c�F�m��@�GoY��'k��R'�u�h	�i�(]|?[Yux��M�SE��]��3�\	����d�Cb`�(�G�����yRv�|��|���X��0@i��o]0V� �=�hw:�E�B�C ���V�Ёt�p.˰�� _�e�i1�_-k�S2q&�o�1��tD�r�9����1`�H�/��_0Yc�ka������M�Gm!�ed���tZ'����`�DQq�����n�L�+U ��)d3Ʈ����B Q�5ya�!�F������v��Bg0$C��/�0�r�C�)Oi���`t��bݫCϞ������<I=(C�NUb�9|%�T��
f��9��MZ>���[�"�4��"{��/�b >ጅjGL�һ�,�Y�$D��[�z���|�B�x�,O$F�UӏE��A�"3�+��Lӯ9:E�V*����Є6ߛ4��.�ٌ�rE�C�yz�М��!�ʁ��Y��D�T,&ϸe�q�׿���
H�����@~5ٕ����T֮�G�lU�`�<C�W��tm����V��ɪ}�#�3�hҺ*&T�m��e�V�1
S -T9�ϗa�;M���W5x%�@uFʬ�K5};���~�N�(M�ƥ[�>ټ]w��Zʗ�0�gw��sq`n�t2Ӥ��Ͼ�,#��ԓ���nQ�С��{���
��(u�@�d�!Q��ߦܙ��=gS���z@R�޲�����KjM8�0X@?�<	��;��)�r����j.k���y�Ȳz�/���?^�&U�Z���e|��/�7���0Ԁ-2m���}��*�XS��Ih9s��<H�F��'y�E��ߦI�p�P�CA�l����q�Iwq�^Mʙ ��a�+���5�"�KI�����ѻK5��br��M���&U��y�����Pp�F��|��ٟ�qɐ���q�C�I���D�� �a�ާ���TdD�˩�om:�I���s5f�u�����S�{��I�G�œU�D��b6�#}�Vv(���R˄G�b�#���O&''��L]�||��}'�8&�d�����r���I('��mkÑ���O7�\�-l߅�_��j,�?�1<�FI�o:h�>z��b	5_7Tihd$���3��ɰWv�%̮̭{WK�2Tf�!}���]"9��98�Ԙ�ö��o���ų�۲	��� ��/�y"��f�狥�?����p#Ѷ��.y�>>����?���ߵf+�1��)mؿ0�б'0�z���O��M�R��D�ǥ�hE��G��i�"6�Vk��RRInr��,є5-8�[3����;'�2��M☐�p�F���^�A>q�J�a̙K��U��\(̣�?�>�}~��0�����{}D�xaěw�'��s�P?�|k��h�K��&��B�]�d�ƈ<d����,�`Ij�xe;5e�����w �$.��?�'�}��:�]#a������P�Fq��Pn��6	�%���fw)�<4GM�Pl��а��q����P��Ư��/�� ����b�}�B4-o�@����M��N�G	�[+C�W�'���w�Z�,ߒ�O ��_�}>(����¤�;�sGlOo�Ŏ��,-�Y4�/�"�3fa��b����%���,�՚�!㦓��b��c,o��۩��f�.�+9B���H��J����b!�מx﯎N��[��ix���r��y_����Sk����GIm�[wt܍���`o���L&9�yґ��*����n��'$�?�I�i`�T�#��j�j�5)o*)/�h.h�H|�?����}%��qd{ f�,����E����f����om6��ρh����>�G��v-܊hc��8L�&_�2~��-���u�5Ht�LZ�
x&��L:(�}r�HXJ��>�*�ez��ο�"�������wl�7���$��e�]��bb��bF��uG,|&�ag�X��C�5����wH��vH�,�;�w���ZCy̨����|�㓎U����%r�j��T]_�J�U�|s&r����	ZJ����[��7F�a�jw��W��1�����8׻�~V��GO��Xs�Yǌ�}�V�ߒe����� .�~��dm�q��j���C�CufM�<C���s��}��j9������u{����E6�3�G��m�w�BTz��6>�_޽6�c��P�Hw�.�9#kR��/���9�B�2C�_��R�|6b��j������x�8�Ն��B;���)�}�o;/ږ��zA�4r�e�c�zA��=^���H�c�z���K�@�.��Vy�5�`���F(��Ċ�d��/m,����=f��_`�6��z������ҍE�ݬNf"�������b��ɘn��w�����:c�i}�4�\h��h��vp�qf��V��X�������]�G@����q)�������e��9&�Z-�rLxC�����k�&Ә�5x�t�~�'>���j���-ᯉg�bI���}'��K4�r
��˦�$�������Ys]�m����0�y��%o�h��LMMM�-��=�R��k�}(���Sf�R�JϳU�4-Ϝi"�t�7D�Ϗ�O^}'UG���F��\?��%��?\3������h-}t0�dʈb{�j��tpuCC�jfwy���י����1�*q�ej�2K-#�Z���x����8;�ݰ��q��fＢl�L/�P	�j����l*�Gf�`t#������qp<� ����E�<�zg�Bk��[܃�?��&��{�g��?PK   W��X�7}b  ]  /   images/c5f41113-5d7c-441f-ad39-f06af9a8b0db.png]��PNG

   IHDR   d   3   ai�   	pHYs  N�  N��"��   tEXtSoftware www.inkscape.org��<  �IDATx��\	��Wq����c�{gfgv��5۬/��)F���("�X�+R!"F�����#Aز�m6���]�w�;;;�s��3����w�����O���.�ݖ�7�]��zU��ޫ�^�]���>D��)wb�d�����p8J�M��x�Q��iH�xڇe�3̣��zI��V��ϝX&��\���U�9��:f��h�P���$X�pbf�!oV�+��
h������i&�j�fJ���Q��0��� �97:�bН%)���#F�w����<�%*�V'��z��fs��Qxg:f	��P
5�����i�Iöi���S�o0y�����)�C�����Q��7�{� 3���p��ӄQ�PG�!�U��;�a:�L��	̡�߻�s2�k�2�	�;�����8�eH�<J�Q�"ux�n�`DC&'��`�0\�`�5ޥ@z�, a_V�i�B�=����e����qd|l������E�{:ZW� ��E��{(Ң{��v!f�?Y�������)wsǌ#��q<?�B�%�*����М��B����ᖫV���qz�O�T���L	���&X��^ӖAS��'φ��u5���˵�^�:nqî$��������ݽ	��fI1�M}o��!�v�8�v ����XN�7���1�<�䲻����%0���ଯ���z�486v�3C3��SC!5��jΡ�)�Gτ�1)o���
�}��Q���Od�b�Nʏo`�)�ߦ�eXm�ؘ�.��ߝ$'��F�%�􌏤t=�����6�`��[	�$t"f@��D�If�ҷ���Й��I������^"WXc,!X%�6M#��(��"b�;+�$ac~�c[rK�J���.��?�u�|h38�X��k�R�f���1ˮ�W�c��^Ni&�X.�*نd�K�,AzYU�λK�D�E�
�'=�$uWI/�F�%�ؕ�`)��� ;Bm���:�t������7#}s���D���Ӥ�]�0���ۚ9ƶ��y��ʙbO�g1a��!�b��o�E��I.K+(�ؠ�P�pV"m�M�M�QOjP��2+o��l�4%@ӯ@_�`3�-�dn�k߇���Ͱj���c��H��drVJr4& �t���	�'�u;������Qlܽd���\T�E��P�D#�9�&"��^�	�6U=a��(ڝ��r�Rdx��!���(�</F4j�%�l�g���G��w��[xn��"�V�n�S���,X��1��V�4p���t�&Bv��P�,a��*	n3� �A�4�{�}���y�m�h�#�����(��wt�&Lj,����,����&��6"�/���4�B�p�:[���#3����Cس�C�?ta
��*Zښ���$��S���mGMM~�h`t|K�q�j/�~�&摜]$�;��gjk��,�p��d����#u����1��Z�;��X+}��� �UD��W��u#��`�ܸ_}C#:;��Leqfp��\�����	~�|���R�>�g%���㖲<�2C4|�8�
�Ģ�R%���l��M�%�]�o��d��	��H��Ko�V�5d`]N���ʩ���P���ġ���IֺX,PZ��2Lw�|����@*�&"9*�P���JR����&L����U�A��ԖN�x�j��`�}�v)U��_P�.]G.WRmҏ9T'���ߔ>G��K�_�Z��TFn�p�o�M��ot|Κ� �t*'F������
�h�Q��ф՚��XM��K�Ee�w��9�7=�$�`0�g���<�BmiV��Ό
���C��C�E ��@3��Bx�0>9O�Ε��Y���qJgrg!�2����2S�o�����ĩ��*��R�X���s?���VI�%$��a���vQ�]�Q�l��W~���tn�qc�[����L$�B���-x�bi���� �����N��l ;щELN/m��%1dc*)���'M-��1��b��084����;�N�q��I�����M��>���<�+�&Hsش��%uLل-�V+GL������XZZ�]w���_����'�p:���[m����xu���ɞ�������Z%�����u��O�63���"�m��������ӆ3���'n;�mm�HҶ�c��<r����|5�UV�|m�k�:9!�M/�gf�h�D[��ر��BKf���dd��%���<v6���r��Ѿ��ؠ�B~L�,���w|�3x��1ڳu��u�p���ٶ��,f
;����Rf��[*����,�y��7�=�N݃sS<��������*�F��jIL_�������S�s�\d���=�C��`�LY��>İ�&sCG�_�닸��G������|wC|��{��lY#������S��u̷��3��1C�]�Cf���&Ƹ���?��]�+9��7<C*��$�.�F2M�By��e��/��LF}��9����s�o?�.4ԇ�9��lr�Y?�啛��ێ��%�%Mՙ._U�,�6�ȯg��c�V|ʕSY�T�������(�JkOkR�07V��夻��V�; Q|�t۠�������(��ne�uy�:K~$�����o�:i	g1�⛿�AW�Mi<p��*a��.F�.�ZBg
z��x�/#\X������W/�POL���tgwCڒ���̹_uy�J3�
.�dc����ئU
۔]�)a'.[�����zJ�y��Sg�w�eqxw�4�//���L�d�t�^S�&u���C�꼁w����l�S�P�:����V���|܃唛�*�Huu��S_bWJ�oL��*��ģ���>�V�8�>O�������n��c��ӆ��9!�}��/h��c�rN��li�E׎f?y�޴�ӋXX\�C,���	��I������D"]�������*��thW� a5ľ�;n^�(#��K87�ώ��:� �O3����������o��_�^o�� �M ��������|��9O�L��_�w|���G߇��>bPZ��q�¤����j2#g���`����� O<����0�����<�����u�a2�����MfO�[ɠ��Z���S�g�3r�~����ŗ.���dp䅳��Ղw�z-j�|ph�iF}�� IG{[�̚���i�v2Y�ֆ09� G��\ՅPЏ=�;��{�M7�G��f^A�sYe�g�o�$����h�S7Y����5!>�|�]b+�6̱Cp�������VM��A�0��3���~�� >����} m��8sn���b��S������8���)L.�֫,���R*�Q��b�:1Ad)N�B�ňo؇G�|ѕU\����)Qao��]�z4�u�"���BLȡ���lC1켨���%��.3g��<Bjk�;���݊���T�V]���ZA�/���Gv�3��n��:ë�'|�$:k�djR�=�����f_�x��uV�RM��5�J;l+N�ˌ��3��y�lۈ���Ɍ`f2sy�����I�5��f����u�)�3���o�&vܵw6�=�p�/z�qg��n�^�sn;��XKj���;*�)֗S�e������Z��՗�Nx�{t�5����U�I�����:�d�{�� �E1�LM��e	6_�s_�.���W�L�h���λ������M*]'՜�����ǃ��O�^��
3!�+��<Fj�g�f�`��p�>��>���y��� ���7ϋ�2���5��͠���o	�xjU�d�����u��� �mwh��O�����+���]�;���j�q�����a"�W�Q�R��g���|a�[l�����L}n!Vv�t���k�z$���i�V$2.��mf��VY��Xd�*_T�\m^�jȞ@�&�~&�����m��28;p�--�����S����h)�yѠ���r�U��y+Icf��qo����=Q�U!�Wބ�ZKl�x���ބ��(b�8��owbp` �@ ���Sr�w���jo%��K5��J���ϊ��nI�
�3rE�kz�c]^��$/��Ey/��y11>�CC��|H�i	~��W���Č�]��юK��_cؐwv��ҒB�z%��.�PЇ��y���������;�W�]C����7�n��KM���'�����;W�0艧^Bm����rs��sϡ��7�r���En.^n��b�K�tPn���U�Ea���M��~�-�ު��iټ����M^�b	�������x\�`Ng+��pb�1�NDԫ�-�e<؁�#���'`��m�\N
��3rH�ʤv�k��H����񤱶��v��&5`Xul�z��Y�`��꟫���G�	&/������tխSG�o����m���6e����>�ۉ��4���G�mү�򂊗Y�)�B��+'Fpwo���W�i<w������߅��Z���3Y�85,������\�wp�.q�O�,b|rA}�v�s��%��oO'��=�L���:����?o��}t�h��؜<.�r�!�n/�i��>,���xF^4��r�Į��]��������s�s��ӄ���j���*F��RG��/Z	���=ޗF�u�^d�"��3gǅ��a|��ߧ�[��b�)�Q���(���y���~^eXXYB��Iĭ�|�`���I:�f��+�����D���-={�/,��cZ2�$lq9A,R{%�J*O3o��f��Nb�I��/�^���ȬH3�V�g
>�OpD���.��0F�%-m��T���r<��Ub�z�-�+���g��$p,�[̀{M�E�2�8'��-l3d�	����)�!7R�]�ɁD|	�ļ ����`bb���sI�K�4�#q!�a�h��[o��))ǁ���U���e5妁�H�F(�L@sx�r["6�Ċ������C,�����KF>���*�y���ޟk�o���22Ɉ�a�R��,]�*r!YD<�}����1��>L�1h,��g��D�dB�1ᮤ� �?GDP�+E��H����Vy���R���6n�yЛE{m\�ۨ�.ڿ$J	��9�連)��@$F] %Ag�eeM"�p���`w��8� �)�j���ql���0v�.��l܏�d������.�f��9ڄ��hJ`;ڄو��&8��S4T���`Rpb��,�֗�ߓ�%I``cZ+�E*M�m��J1ֳ�2�8��͕��fH�̢�;�Z�#����q�1b�	qdP�:�!W�Ys�S��80�S6��r�KĔ�Vua.+$�n�@H����J�S�7�'PD�`�DtuH��ƣ>�R�C��� �0��5��T.�х�!�R�M���c1�<u�nn=�Q(2���fB��pq8𘄧AL��Q|�.��7$<��R��M��� a��z�����k�۩�����o�|����l�WgZ�眛�єV����2¤�-�7KOc�.Y�rT9&�N��s�F�2��2��)<p�N��%?�1$��'�T�	�Wc&�N⡗k�-ZoΉ�o#�/�D@�0�����^��-3��p�R�f8�U�9�{_{�F��)���а�9+���p���b`+���ٰ�&�1��ud��S�"�<�0G,�MJt"���@~��^b����jl��J%C>C�����,TȠN�����D��χ�s(��[+�i�d�T���OPqY0V;cKLF��rr�鱁�2�$��	_y���-��,��c*���\PS����G��̡��0�ϯ΅����Ϗ��ݹ�h@چ�G<��S6��YqK@a�5�(1��ӢT��d���OBE`�G���Ǳ!�ɏ,6r���]f��$�ӎ���3D7s�2���G\k%�(G\sav���}������k�f�6����0�;Ov))1�x@���۰:�J���a�r�yC!϶��b�hk �dG���Nd֢ޑ�X*���^�.kE�c��ޱ�d|�g�D�c)ZQ�8��4{,�������L�����a#8�}�t�?��q�d�    IEND�B`�PK   ��Xx*�X  S  /   images/f4d2e4ba-8b5e-4c52-bc1f-19feb473bfd1.pngS��PNG

   IHDR   d   p   ���   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��]yp�e����;�NH�A �0
r@��Q�Y�rtX�ݲԝ�Úuժqg�f��cj�vV�r`Ww���U\t� (�B$�s_�������_h��:�N�n~�[!ݝ�����������fD���:���򿿕�+i=>o���,틿�Q�On�$҈8n�N�u�4�����*�٣-gT	q�\�ӥ�x[Le��Ț����	u�j0�H�C|=�H��9��p�*!w�qz�A̚5�ן\���T�={O���~��3g�nw@�d,//������,#!�$�a���[����/����j�/��^7x�����ƶ���
���/^tKs-[���b�4���>r�d25��mۄ���4x�#���9�}h8B,ҶJ�)|�����k����V$�)^X��*���(���]iwI��P0B(�+�n����1�?�g��)z���W�m�"��k�����ɸc�8�$����O��.�/0�hc=<cMR��j|	I�~�C����1�oQ�h���ץ��ג3`	��ͅ�h�N�>p�� �Á��FՂ�
���]���0zb4�K��l���_�+V ??_�>���	��ׇS�Na�Ν8v��G9�Ԕ�sdߓ�J����x衇p�UWappN��a�� ���3f`ǎ����>JM�IBV�}�d2�P_H�C蠖p���y�����_�昫�ڞ�+WbΜ9Aɠ�$q��& �Ho��ǂP����7��v�������s���b�^{����@TG2��Ѐ��fuQ��6������'+�~��������`��V�U�;//O��|mܸqX�h>��À߯K����QXX��I����O>AKK�e���,\�7�|�
~,>��f_>��c�o��)++����ڵk���7ɚ>}z���9�U���n��͛U�P^^�k��{��Ņ�g:;;��T>�-�I!x��p��5���ϫ�	Z��?�\�����W�޿�4m999���%�������n<��38s�֭[�ŋ#==]�,����곏=�&N����dǢ��_MB��$⦛nBII	�oߎ����>�	����G��i�B�wH	g�i�q�-�`���JP6�h ���_~Y	ǎ%c2IK��{�)2��ƍ7j��#h����\��o�����	�vPv�ޭ�Wee��b2�}�ހ�#G���ٳ��t������o��lذA���b�@���!��G���q��	�y655�^P|�W���-##CiD |��wʦ&��'��<QK-�=FU����*B|���|٦Cg���T��|������������姟~���
̟?'O����Ģ�C�5�ߩ�r'�b���h�؆��o_s!��H@�KO�~���S�����)S���&P(�蠙e�����eث-�h���P���25�tI�ܹs�2a��oБ��D���G,��BV��z�شiSH��K	*_��^ms�i��+�!���3|���*t%l������u=���Q�u�]غud�SqS�nu���wyU�$3�"���,Zg��@'�5���)���+�� ��=u�T�{�x���G4�,Y���P�B�[�5k�(g�e�v�S��%�@8�F4C��q�V䵴"���Y������!�7-�9Yh�<������̡�
�j7W&�����+?X&�@3�>�jV� &b���p5�k:��Ç����0F��EEE곡��lj�E��҆s�kmG�����!���wh�h[Fo/�[Z0�����ج�/-��ɑ�1��[j�S��wNP:p��f��ND��8�cf�M,�%m��g83(d8>�f&E��r��g��խ�nrIS&��(u{7|@3���{_��=�_��_lFq�Etf�DM�$ԖOB��fS���I-�
75F�7C[-f��[���
�ڠ�Bl�FRj���Һz�<v��.�I���S�h�QL�� _Z���4x��H�ϸEW[��Mp
.ɮI��O�zz1��{�՝���+� Z���A[8���&�X����#���]&1O�}����՟S�!ES��`�4��4������<vN����W�!S1G!͜_ ��RE�`SN�z�E͑�#��d��il��f�!�kt�nb���ҐH��+�~�7��&�Z�ɄAl�0�F�ė���gC�����pj�U���S���?b��f���6�#El�g`k����W�U S����J��B#�?�4�Ɋ�Ӱ@[+,bR�Ԉ�]�����g��_�e%�頵.n1k����cU��5mb��ه}�碱�0�$��(2�_�����:5�L��,�to������>�`� dx��e���7\���+��dB,��_/�'��MS�B��k�+Ͱ:=�'�*.6z���ϰ�� !���B&MJ�B���\���qQ#%�4�-�R��΅�3RE����ɠs�-���^��x�CJ&G(�(���T*GopE~� �al;�j�r�.��V2bom,M�P��Q�}� ֈ)!$������_"���Ŧؓ�a����DEf��26JbZ;�<�+!4��_�$e3����p ��5�/h拲{~)kca�Zj���q0Č��)�k$S�m@_o|��@(KG;`�SD�J��%q����]C��=(�����ޒ�D C�6I2�T8LY������r�����ĄvlB�9�d>����u�DA�(��(j"��)�OVL����]CLb�'4��,�k���9�� T���EK(3|͔��uB���6�::�֏�ӝ�ڡ��QFk�G���)֖kS�(�E\5�3,_�rn�g��ݘ(�4���9;>�#���y����BG8N=?�c��{$�v�s8�$	b�zt� }h��dw�����٭�L�bǜ	M�=]��^B�b��'�g9싓��$&��"ڐ*�mH��
M�T����U�-���}��7ʏ�G]CR���?�$7��Y4�^H)L��>�/=��ɭ!�[uܗLV��!��seZ2wn�Zb�lK�5�#�}��N`��O�SD�FG/\�{]~g_�p}�M};���<h���0(h��č�۳��{SӪp��$��GL�$�)��w�(|�' ��!�����p�9ef�I����e�:�.�K��r��m'�QC��6N� ��;������N�ݻL���Mp��D}�7��H�N���"Ul1,�P�D�
����sb�Rd2q��RS�/����?�.�vtdg�:���N������ې��y��������Ď�l�S�ɋA�%Z���I��TGMf�:������-2�3D3�0�G"%�}q�9dv���ǧ��ssUU���$�������w�bV}����+!�?���j�����3�dw9a�-H,P;ZE�����(Oˀ�jU}0��/ml�p�<�-����v�c̔Y�U�넜���͢{5aJ�PCO(V}��l�rf�+)Bŉ��u�c�5�S_���a.$��2��3�d�fee�m�A��� bB��Gd�Ք��Z}s�6�p����/32U��0���%2��41��D�Se���?�ۀ�0>F�[��{zP�;��tWJ�;גw�ť�������e�h����&F\;�j	�髞Y��U�2� {[�x���F�4#�S�A8/�]d����,k���钝���ф���ˎ��P��M1�L=n�N��P�{{�.+�QDl�h(C׬�U��2_9uQzN$!4D5��ʙ����*�������=��k!%WB́�'I�ZE���k�Ind���	]2�J�rF����E\��w�����}�yI)��9��b���ݍ{2�1�d� ����왟�[�Y���&y�"䬭��S������Q��JC�,��������?	��Q��!e}Z:[,�U�_[ۋ�J&��Qu�s^ILӍӮ@�u��"I`4�F�B�í���٢X�� �2���,:���ĞWZp3�y�ݣ�UH�I��kT�;�$�P����<���+*`Y�M6[\�č�S����\|�t*��~��$ep��>*?��,W"��hFA4$Ù3�]��o�,1���R�B��[��B'>w.2�4gf�2RC4��Z�{�B�ε�o�ӱ���Ŝ�ɀ}�p`�����L��y���:���+5���q����zhp ��g/K��I��mr�y+V e�bt�0M�1B��T��O�Z����
��Å8P]�?�/��A �"�<����јq�3K~O����$���Y>���;����\|�W~�����f5ܥ�'D�p���9j�b+Z=t���X���� ��'���-��W��.��iS��P5;����d��������d�����H�g�ڠ
�p��q�I�P^Y	ی鞛�IP��f��a1L6�����
�I�	�N`ͨ/��R�BgYq^���X�h�ҥ�\Q�GW(m���e��b�<L;q�Ǐ���ڄx�$�6C�L��u��s?�|.Ed�M���9�a+/��;p�޴�kr�4,���O�{�
*��e��.KE�L����o��4�$���Nն]�z5n����E���EiCa>LE�Q�x!����jh@˹sh���-��:�[U�y�n��lM�Z�YT�ĉ��� �[ ��	���3���>����
Xǘ�"���ρH���p����[x��"���qf����EY��GY��$�]83F�-(S��79��XZ����,��J?l,���~�]��h��u���X+;�e�U��U�9�,��R�,E��Ť�mۦ�.��@f;b�p��߿_��
jw�}7JKK����@�Jفw�yGi�h�.�ej���t_�h�:�%��L�>��7�T}a�\]D�́��(��h`�'��bU�P�R�q�j�O�HyQ`���1���6¬�
��<#d׮]��;OF`%=���}��
�����CD4D+�___�����Ԏ�cX�
�$��Y2�꿳ߔ���vh�L����KO�>���xek
������O�h�E!MQp��S�d��N�);���%�� �d��s{)�Z����N=��C�40��icltr�H��&�v���k�<މ�X�r�#=z?b�0�	�|Áɢ^�De��@�2��L!���:��_�>@�){�u�5�o�5"b���+���E�����xTe����~�˱�V+|B�C#�1C<�/���������BǊcJA鐋�>#�	�81gIƳC4hy�ٳgUI���QX8���"����>�_|Qe����y�$���t6_��?��:X��E00;����V}����]B��0��~��~^�'p}j߾}�DO
�]���W���Z�Je��L�����drᔫ�<�Kp�`\*�*Oe�ʏ��c�w��K73sV��gT;���΋S����׹�Ŭ��Q˒�o�}a�N���:u2�Fb<6��Y[���s� ��!�,h楝Nb����C&}���ؠ���Sch��C�;�5�	㺞o�폠�p�lǎظq��
j�������cG���믇�I�c��M�܈�� fg��6��0,��<j���W_.{��l��Śg�>��g��5+.��*��dcc���^� �m��G�=���?x���*nLi;�c��H����'�_BRܸD�.~�;N�Gi������7�C�f�!�i��}!P��R�`�M��/ꅽ��p�sC4�4<N����	M��I�G?���p���KsH���p�������7�嗿0N�=sfw{{{#<7���U����ye���q���]�O�!��9�|����`���K��P^�f�?I�D���V믶����f/�4k.���/~񉄩��ߗ������y����#G�*K�G�\��7D��k��-B�I�_�w������~Î;R7n������&��D���^{g��;�`0��>/�b����q}���+��F����#$��BE0`zR�    IEND�B`�PK   ��X%P��  �     jsons/user_defined.json�X�n�8��Ϧ��%oE�]ۦEnX`�-֑\InP��IIӆ�Cg��X4OE�!����n�}Y���|ӆ�����/�CӖu�/	���Om��=�s\����>�;<�]�����J	�]х�����o�.4U�fu��]��U;�\!��#t�&,�%��k:�`�AL񀬣1n0f�F����5�W�8��t=�*����"^���QL�':H��r]]�{����%'"'�0$�r�sQ�A�"�B[���K7�Ux[�f��+����
w�麬�T���ͫ��QٮWŗ�zI���1���Է�3Hz�7B�)�T��z�O�r؟M?�n�>��r#T���,���b�(�W���x�!ѫ~�+<���Np6�+6	�U����G��4��#������,A=:0G碟�It���q�f��It����lt2�.t=dF(��~8��t3�K��>MI��<��lN��1	oRx2��lN�<I�JF���v1�K�j��5�d3���4~*Z2�VJ�͞�ӳ� �n�p)�9G�J��1C|�f>�;06 U/�zɴ�ja��r8�]�vT�T�l�g8�<�T�|�',���TâG�D�|�HE,��+e������jX����ߥa�jX��D��`�ś�،; 2?Cb���xd��� [4L� ���@MH5L�",����"&l8d���ɟ�R�Qƒ��lG�-W�cL�u���[n�AɊ�|%J�����ܖ���0����t�`i`��o�u������~m?Z�����j�f��✃��=���{'c�pXJ���qb(*�H.xм��u�%�Vw��x����`��̋i�d�A�0S��1X�H9C.�IQ�M
�#C�-
���_;��TH����R��JО1��d�4���So�}�|�	߮*����.�	�g���2�mySv�����uw�Q�h��"�0��D�`́�E_^JSx�S+9"�>��@F�Ɯڂ+^��{���4>Õ�pJ@�c��O) �P'�f)9X�ݜ��C[�<��3?~����?�-���B+�A{(*D#N1C��"6�YMU����ֶ]5$e�M{m7]S���h���*��t�Ł�SVcP��X0�\��[l)@~��~M%g5C�K�8���0�T����AZ�T�ҭ_~���p���%�R�K��s~`h��K߁/� B�g��G��)ucK8�S;�`��N��� �l�g����;j;Ƈ��{��Y��Xm*��!h�d�5Xtwϱ���}uJ�����e[�U�6քO�!�p����b�&��4��.� ��6�O��C5����m����a�8�#*{�B1=��TK��֯�ePp�y��4�͎R>�@��
*�$@#�6�H�9Wدj��������+$�j����R�Xɜ	�W�˯� PK
   ��X�zG��  �K                  cirkitFile.jsonPK
   ��X��.P9  4  /               images/3f03cad7-594e-4892-9bc7-779b63c9e608.pngPK
   ��X�"{Q�? �f /             �.  images/4321cb83-9d65-4877-9350-be2835182319.pngPK
   ���X�ة� � /             �n images/4cb229e9-cddc-4c52-860a-b86ee61c7037.pngPK
   ��X>6YYJ �r /             ͈ images/54ec96e0-e6c8-4747-b5e8-2cd896730fff.pngPK
   W��X8�w���  ��  /             8� images/805fb750-7b5b-4a1e-90f5-2022d18e6d35.pngPK
   ,��X�u�Q�"  &  /             �� images/87392e8d-b818-4203-815b-f0983b827fd2.pngPK
   ���X��/F��  ��  /             �� images/906ef243-ce1b-4f5e-9eb4-92ebaa7c38d8.pngPK
   ,��X5��<O  g  /             �� images/c0642b64-198f-4d8a-96f5-22ba47d3499f.pngPK
   W��X�7}b  ]  /             H� images/c5f41113-5d7c-441f-ad39-f06af9a8b0db.pngPK
   ��Xx*�X  S  /             �� images/f4d2e4ba-8b5e-4c52-bc1f-19feb473bfd1.pngPK
   ��X%P��  �               � jsons/user_defined.jsonPK      $  �
   